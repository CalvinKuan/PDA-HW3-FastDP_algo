VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LAYER LEF58_CORNERSPACING STRING ;
END PROPERTYDEFINITIONS

CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.0005 ;
USEMINSPACING OBS ON ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.0115 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.50
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.10        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.28        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.50        0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.06 ENDOFLINE 0.06 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.014 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  AREA 0.017 ;
  MINWIDTH 0.05 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  AREA 0.025 ;
  MINWIDTH 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.15 ;
  WIDTH 0.10 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  AREA 0.052 ;
  MINWIDTH 0.10 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA12_PG
    LAYER Metal1 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via1 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA12_PG

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_E DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_E

VIA VIA23_1ST_W DEFAULT 
    LAYER Metal2 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_W

VIA VIA23_PG
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via2 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA23_PG

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_N DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_N

VIA VIA34_1ST_S DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_S

VIA VIA34_PG
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via3 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA34_PG

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C

VIA VIA45_PG
    LAYER Metal4 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
    LAYER Via4 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
END VIA45_PG

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA56_PG
    LAYER Metal5 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
    LAYER Via5 ;
        RECT -0.150000 -0.150000 -0.100000 -0.100000 ;
        RECT -0.150000 0.100000 -0.100000 0.150000 ;
        RECT 0.100000 0.100000 0.150000 0.150000 ;
        RECT 0.100000 -0.150000 0.150000 -0.100000 ;
    LAYER Metal6 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
END VIA56_PG

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA6_0_HV

VIA VIA67_PG
    LAYER Metal6 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via6 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA67_PG

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
END VIA7_0_VH

VIA VIA78_PG
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via7 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal8 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA78_PG

VIA VIA8_0_HV DEFAULT 
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
    LAYER Via8 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal9 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
END VIA8_0_HV

VIA VIA12_2C_W DEFAULT
    LAYER Metal1 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA12_2C_W

VIA VIA12_2C_CH DEFAULT
    LAYER Metal1 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via1 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA12_2C_CH

VIA VIA12_2C_E DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via1 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA12_2C_E

VIA VIA12_2C_S DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA12_2C_S

VIA VIA12_2C_CV DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via1 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA12_2C_CV

VIA VIA12_2C_N DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via1 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA12_2C_N

VIA VIA23_2C_W DEFAULT
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA23_2C_W

VIA VIA23_2C_CH DEFAULT
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via2 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA23_2C_CH

VIA VIA23_2C_E DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via2 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA23_2C_E

VIA VIA23_2C_S DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA23_2C_S

VIA VIA23_2C_CV DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via2 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA23_2C_CV

VIA VIA23_2C_N DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via2 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA23_2C_N

VIA VIA34_2C_W DEFAULT
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA34_2C_W

VIA VIA34_2C_CH DEFAULT
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via3 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA34_2C_CH

VIA VIA34_2C_E DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via3 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA34_2C_E

VIA VIA34_2C_S DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA34_2C_S

VIA VIA34_2C_CV DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via3 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA34_2C_CV

VIA VIA34_2C_N DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via3 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA34_2C_N

VIA VIA45_2C_W DEFAULT
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA45_2C_W

VIA VIA45_2C_CH DEFAULT
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via4 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA45_2C_CH

VIA VIA45_2C_E DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via4 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA45_2C_E

VIA VIA45_2C_S DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA45_2C_S

VIA VIA45_2C_CV DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via4 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA45_2C_CV

VIA VIA45_2C_N DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via4 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA45_2C_N

VIA VIA56_2C_W DEFAULT
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA56_2C_W

VIA VIA56_2C_CH DEFAULT
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via5 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal6 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA56_2C_CH

VIA VIA56_2C_E DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via5 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA56_2C_E

VIA VIA56_2C_S DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA56_2C_S

VIA VIA56_2C_CV DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via5 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA56_2C_CV

VIA VIA56_2C_N DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via5 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA56_2C_N

VIA VIA67_2C_W DEFAULT
    LAYER Metal6 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
END VIA67_2C_W

VIA VIA67_2C_CH DEFAULT
    LAYER Metal6 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
    LAYER Via6 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
END VIA67_2C_CH

VIA VIA67_2C_E DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
    LAYER Via6 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
END VIA67_2C_E

VIA VIA67_2C_S DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
END VIA67_2C_S

VIA VIA67_2C_CV DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
    LAYER Via6 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
END VIA67_2C_CV

VIA VIA67_2C_N DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
    LAYER Via6 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
END VIA67_2C_N

VIA VIA78_2C_W DEFAULT
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
END VIA78_2C_W

VIA VIA78_2C_CH DEFAULT
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
    LAYER Via7 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
END VIA78_2C_CH

VIA VIA78_2C_E DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
    LAYER Via7 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
END VIA78_2C_E

VIA VIA78_2C_S DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
END VIA78_2C_S

VIA VIA78_2C_CV DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
    LAYER Via7 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
END VIA78_2C_CV

VIA VIA78_2C_N DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
    LAYER Via7 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
END VIA78_2C_N

VIARULE M4_M3 GENERATE DEFAULT
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
END M4_M3

VIARULE M5_M4 GENERATE DEFAULT
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
END M5_M4

VIARULE M6_M5 GENERATE DEFAULT
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
END M6_M5

VIARULE M7_M6 GENERATE DEFAULT
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
END M7_M6

VIARULE M8_M7 GENERATE DEFAULT
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
END M8_M7

SITE CoreSite
  CLASS CORE ;
  SIZE 0.1 BY 1.2 ;
END CoreSite

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.010 BY 23.5000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 23.5000 BY 23.5000 ;
END corner

MACRO XOR2X2
  CLASS CORE ;
  FOREIGN XOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.685 0.171 1.748 0.998 ;
      RECT 1.655 0.171 1.685 0.395 ;
      RECT 1.655 0.693 1.685 0.998 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.368 0.564 0.461 0.694 ;
      RECT 0.326 0.639 0.368 0.694 ;
      RECT 0.263 0.639 0.326 0.763 ;
      RECT 0.239 0.706 0.263 0.763 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.869 0.499 0.931 0.585 ;
      RECT 0.686 0.530 0.869 0.585 ;
      RECT 0.637 0.530 0.686 0.630 ;
      RECT 0.574 0.454 0.637 0.630 ;
      RECT 0.229 0.454 0.574 0.508 ;
      RECT 0.166 0.454 0.229 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.533 -0.080 1.800 0.080 ;
      RECT 1.440 -0.080 1.533 0.122 ;
      RECT 0.720 -0.080 1.440 0.080 ;
      RECT 0.627 -0.080 0.720 0.122 ;
      RECT 0.305 -0.080 0.627 0.080 ;
      RECT 0.213 -0.080 0.305 0.122 ;
      RECT 0.000 -0.080 0.213 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.530 1.120 1.800 1.280 ;
      RECT 1.437 1.078 1.530 1.280 ;
      RECT 0.698 1.120 1.437 1.280 ;
      RECT 0.605 0.905 0.698 1.280 ;
      RECT 0.305 1.120 0.605 1.280 ;
      RECT 0.213 0.905 0.305 1.280 ;
      RECT 0.000 1.120 0.213 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.583 0.473 1.621 0.558 ;
      RECT 1.520 0.212 1.583 0.558 ;
      RECT 1.182 0.212 1.520 0.267 ;
      RECT 1.376 0.520 1.439 0.994 ;
      RECT 0.895 0.939 1.376 0.994 ;
      RECT 1.245 0.336 1.308 0.802 ;
      RECT 1.120 0.212 1.182 0.838 ;
      RECT 1.015 0.212 1.120 0.293 ;
      RECT 1.091 0.783 1.120 0.838 ;
      RECT 0.998 0.783 1.091 0.864 ;
      RECT 0.994 0.368 1.057 0.708 ;
      RECT 0.946 0.368 0.994 0.423 ;
      RECT 0.895 0.654 0.994 0.708 ;
      RECT 0.911 0.206 0.946 0.423 ;
      RECT 0.884 0.163 0.911 0.423 ;
      RECT 0.832 0.654 0.895 0.994 ;
      RECT 0.818 0.163 0.884 0.261 ;
      RECT 0.802 0.717 0.832 0.940 ;
      RECT 0.513 0.206 0.818 0.261 ;
      RECT 0.717 0.319 0.810 0.400 ;
      RECT 0.502 0.765 0.802 0.820 ;
      RECT 0.142 0.332 0.717 0.387 ;
      RECT 0.420 0.193 0.513 0.274 ;
      RECT 0.439 0.765 0.502 0.905 ;
      RECT 0.409 0.824 0.439 0.905 ;
      RECT 0.104 0.281 0.142 0.387 ;
      RECT 0.104 0.683 0.142 0.764 ;
      RECT 0.104 0.950 0.138 1.031 ;
      RECT 0.041 0.281 0.104 1.031 ;
  END
END XOR2X2

MACRO XNOR2X2
  CLASS CORE ;
  FOREIGN XNOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.948 0.171 1.950 0.395 ;
      RECT 1.884 0.171 1.948 0.998 ;
      RECT 1.857 0.171 1.884 0.395 ;
      RECT 1.854 0.693 1.884 0.998 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.490 0.564 0.521 0.645 ;
      RECT 0.427 0.564 0.490 0.694 ;
      RECT 0.402 0.627 0.427 0.694 ;
      RECT 0.329 0.639 0.402 0.694 ;
      RECT 0.266 0.639 0.329 0.763 ;
      RECT 0.241 0.706 0.266 0.763 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.059 0.468 1.123 0.585 ;
      RECT 0.875 0.530 1.059 0.585 ;
      RECT 0.811 0.530 0.875 0.630 ;
      RECT 0.668 0.575 0.811 0.630 ;
      RECT 0.647 0.573 0.668 0.630 ;
      RECT 0.584 0.454 0.647 0.630 ;
      RECT 0.231 0.454 0.584 0.508 ;
      RECT 0.168 0.454 0.231 0.555 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.741 -0.080 2.000 0.080 ;
      RECT 1.647 -0.080 1.741 0.122 ;
      RECT 0.810 -0.080 1.647 0.080 ;
      RECT 0.716 -0.080 0.810 0.122 ;
      RECT 0.386 -0.080 0.716 0.080 ;
      RECT 0.292 -0.080 0.386 0.122 ;
      RECT 0.000 -0.080 0.292 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.727 1.120 2.000 1.280 ;
      RECT 1.634 1.078 1.727 1.280 ;
      RECT 0.788 1.120 1.634 1.280 ;
      RECT 0.694 0.905 0.788 1.280 ;
      RECT 0.380 1.120 0.694 1.280 ;
      RECT 0.287 0.905 0.380 1.280 ;
      RECT 0.000 1.120 0.287 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.781 0.471 1.820 0.558 ;
      RECT 1.718 0.196 1.781 0.558 ;
      RECT 1.376 0.196 1.718 0.251 ;
      RECT 1.572 0.520 1.635 0.994 ;
      RECT 1.022 0.939 1.572 0.994 ;
      RECT 1.439 0.306 1.503 0.802 ;
      RECT 1.313 0.196 1.376 0.838 ;
      RECT 1.207 0.196 1.313 0.302 ;
      RECT 1.284 0.783 1.313 0.838 ;
      RECT 1.190 0.783 1.284 0.864 ;
      RECT 1.186 0.357 1.249 0.708 ;
      RECT 1.087 0.357 1.186 0.412 ;
      RECT 1.022 0.654 1.186 0.708 ;
      RECT 1.023 0.199 1.087 0.412 ;
      RECT 0.601 0.199 1.023 0.254 ;
      RECT 0.959 0.654 1.022 0.994 ;
      RECT 0.927 0.717 0.959 0.940 ;
      RECT 0.862 0.308 0.956 0.389 ;
      RECT 0.590 0.765 0.927 0.820 ;
      RECT 0.143 0.321 0.862 0.376 ;
      RECT 0.507 0.186 0.601 0.267 ;
      RECT 0.526 0.765 0.590 0.905 ;
      RECT 0.496 0.824 0.526 0.905 ;
      RECT 0.105 0.281 0.143 0.376 ;
      RECT 0.105 0.683 0.143 0.764 ;
      RECT 0.105 0.950 0.139 1.031 ;
      RECT 0.041 0.281 0.105 1.031 ;
  END
END XNOR2X2

MACRO SEDFFTRX2
  CLASS CORE ;
  FOREIGN SEDFFTRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.697 0.150 0.838 0.258 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.379 0.514 0.488 0.633 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.260 0.356 0.293 0.494 ;
      RECT 0.212 0.343 0.260 0.494 ;
      RECT 0.170 0.343 0.212 0.424 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 6.561 0.573 6.593 0.627 ;
      RECT 6.557 0.346 6.572 0.439 ;
      RECT 6.557 0.573 6.561 0.737 ;
      RECT 6.496 0.346 6.557 0.737 ;
      RECT 6.482 0.346 6.496 0.427 ;
      RECT 6.471 0.656 6.496 0.737 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 6.920 0.306 6.943 0.361 ;
      RECT 6.901 0.306 6.920 0.724 ;
      RECT 6.859 0.306 6.901 0.737 ;
      RECT 6.821 0.346 6.859 0.427 ;
      RECT 6.810 0.656 6.859 0.737 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.128 0.433 2.241 0.550 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.457 0.439 1.624 0.524 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 3.208 0.439 3.443 0.494 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.741 -0.080 7.000 0.080 ;
      RECT 6.651 -0.080 6.741 0.258 ;
      RECT 6.142 -0.080 6.651 0.080 ;
      RECT 6.052 -0.080 6.142 0.122 ;
      RECT 5.404 -0.080 6.052 0.080 ;
      RECT 5.398 -0.080 5.404 0.118 ;
      RECT 5.149 -0.080 5.398 0.199 ;
      RECT 5.144 -0.080 5.149 0.118 ;
      RECT 4.457 -0.080 5.144 0.080 ;
      RECT 4.367 -0.080 4.457 0.274 ;
      RECT 3.739 -0.080 4.367 0.080 ;
      RECT 3.648 -0.080 3.739 0.335 ;
      RECT 3.377 -0.080 3.648 0.080 ;
      RECT 3.287 -0.080 3.377 0.122 ;
      RECT 2.345 -0.080 3.287 0.080 ;
      RECT 2.255 -0.080 2.345 0.245 ;
      RECT 1.571 -0.080 2.255 0.080 ;
      RECT 1.481 -0.080 1.571 0.122 ;
      RECT 0.609 -0.080 1.481 0.080 ;
      RECT 0.518 -0.080 0.609 0.197 ;
      RECT 0.162 -0.080 0.518 0.080 ;
      RECT 0.072 -0.080 0.162 0.122 ;
      RECT 0.000 -0.080 0.072 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.731 1.120 7.000 1.280 ;
      RECT 6.641 0.971 6.731 1.280 ;
      RECT 5.953 1.120 6.641 1.280 ;
      RECT 5.953 0.863 6.022 0.914 ;
      RECT 5.841 0.863 5.953 1.280 ;
      RECT 5.772 0.863 5.841 0.914 ;
      RECT 4.987 1.120 5.841 1.280 ;
      RECT 4.897 1.078 4.987 1.280 ;
      RECT 4.413 1.120 4.897 1.280 ;
      RECT 4.164 1.078 4.413 1.280 ;
      RECT 3.371 1.120 4.164 1.280 ;
      RECT 3.281 1.008 3.371 1.280 ;
      RECT 2.317 1.120 3.281 1.280 ;
      RECT 2.227 1.008 2.317 1.280 ;
      RECT 1.556 1.120 2.227 1.280 ;
      RECT 1.466 1.008 1.556 1.280 ;
      RECT 0.488 1.120 1.466 1.280 ;
      RECT 0.398 1.078 0.488 1.280 ;
      RECT 0.000 1.120 0.398 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.737 0.505 6.798 0.592 ;
      RECT 6.735 0.537 6.737 0.592 ;
      RECT 6.674 0.537 6.735 0.887 ;
      RECT 6.338 0.832 6.674 0.887 ;
      RECT 6.338 0.162 6.346 0.386 ;
      RECT 6.277 0.162 6.338 0.887 ;
      RECT 6.256 0.162 6.277 0.386 ;
      RECT 6.243 0.699 6.277 0.887 ;
      RECT 6.153 0.699 6.243 0.952 ;
      RECT 6.202 0.464 6.216 0.545 ;
      RECT 6.187 0.458 6.202 0.551 ;
      RECT 6.126 0.282 6.187 0.630 ;
      RECT 5.607 0.699 6.153 0.754 ;
      RECT 5.778 0.282 6.126 0.337 ;
      RECT 5.485 0.575 6.126 0.630 ;
      RECT 5.859 0.419 5.873 0.500 ;
      RECT 5.783 0.419 5.859 0.506 ;
      RECT 5.348 0.451 5.783 0.506 ;
      RECT 5.687 0.269 5.778 0.350 ;
      RECT 5.546 0.699 5.607 0.994 ;
      RECT 3.769 0.939 5.546 0.994 ;
      RECT 5.424 0.575 5.485 0.817 ;
      RECT 5.221 0.327 5.408 0.382 ;
      RECT 5.287 0.451 5.348 0.870 ;
      RECT 3.902 0.815 5.287 0.870 ;
      RECT 5.160 0.327 5.221 0.740 ;
      RECT 5.038 0.483 5.099 0.746 ;
      RECT 4.619 0.692 5.038 0.746 ;
      RECT 4.775 0.231 4.860 0.312 ;
      RECT 4.770 0.231 4.775 0.623 ;
      RECT 4.714 0.244 4.770 0.623 ;
      RECT 4.709 0.244 4.714 0.460 ;
      RECT 4.684 0.568 4.714 0.623 ;
      RECT 4.695 0.379 4.709 0.460 ;
      RECT 4.619 0.221 4.648 0.302 ;
      RECT 4.558 0.221 4.619 0.746 ;
      RECT 4.477 0.660 4.558 0.740 ;
      RECT 4.407 0.349 4.497 0.430 ;
      RECT 4.276 0.673 4.477 0.727 ;
      RECT 4.107 0.362 4.407 0.417 ;
      RECT 4.274 0.543 4.276 0.727 ;
      RECT 4.215 0.517 4.274 0.727 ;
      RECT 4.184 0.517 4.215 0.598 ;
      RECT 4.046 0.192 4.107 0.596 ;
      RECT 4.004 0.192 4.046 0.246 ;
      RECT 3.861 0.542 4.046 0.596 ;
      RECT 3.866 0.301 3.956 0.382 ;
      RECT 3.841 0.737 3.902 0.870 ;
      RECT 3.862 0.327 3.866 0.382 ;
      RECT 3.801 0.327 3.862 0.485 ;
      RECT 3.800 0.542 3.861 0.679 ;
      RECT 3.739 0.737 3.841 0.792 ;
      RECT 3.739 0.430 3.801 0.485 ;
      RECT 3.708 0.861 3.769 0.994 ;
      RECT 3.678 0.430 3.739 0.792 ;
      RECT 3.615 0.861 3.708 0.915 ;
      RECT 3.102 0.611 3.678 0.665 ;
      RECT 3.493 0.985 3.629 1.039 ;
      RECT 3.554 0.735 3.615 0.915 ;
      RECT 2.946 0.735 3.554 0.789 ;
      RECT 3.432 0.883 3.493 1.039 ;
      RECT 0.960 0.883 3.432 0.938 ;
      RECT 3.102 0.257 3.171 0.338 ;
      RECT 3.081 0.257 3.102 0.665 ;
      RECT 3.041 0.270 3.081 0.665 ;
      RECT 2.914 0.645 2.946 0.789 ;
      RECT 2.914 0.271 2.937 0.352 ;
      RECT 2.853 0.271 2.914 0.789 ;
      RECT 2.846 0.271 2.853 0.352 ;
      RECT 2.742 0.645 2.755 0.726 ;
      RECT 2.742 0.271 2.746 0.352 ;
      RECT 2.726 0.271 2.742 0.726 ;
      RECT 2.681 0.271 2.726 0.789 ;
      RECT 2.655 0.271 2.681 0.352 ;
      RECT 2.665 0.645 2.681 0.789 ;
      RECT 1.922 0.735 2.665 0.789 ;
      RECT 2.544 0.456 2.585 0.543 ;
      RECT 2.544 0.279 2.559 0.360 ;
      RECT 2.483 0.279 2.544 0.665 ;
      RECT 2.469 0.279 2.483 0.360 ;
      RECT 2.427 0.611 2.483 0.665 ;
      RECT 2.362 0.468 2.421 0.523 ;
      RECT 2.302 0.468 2.362 0.665 ;
      RECT 2.047 0.611 2.302 0.665 ;
      RECT 2.047 0.293 2.132 0.374 ;
      RECT 2.042 0.293 2.047 0.665 ;
      RECT 1.986 0.306 2.042 0.665 ;
      RECT 1.869 0.267 1.922 0.789 ;
      RECT 1.861 0.267 1.869 0.829 ;
      RECT 1.808 0.640 1.861 0.829 ;
      RECT 1.147 0.774 1.808 0.829 ;
      RECT 1.685 0.269 1.746 0.680 ;
      RECT 1.656 0.269 1.685 0.324 ;
      RECT 1.617 0.625 1.685 0.680 ;
      RECT 1.322 0.260 1.384 0.340 ;
      RECT 0.622 0.993 1.364 1.048 ;
      RECT 1.322 0.639 1.355 0.694 ;
      RECT 1.294 0.260 1.322 0.694 ;
      RECT 1.261 0.273 1.294 0.694 ;
      RECT 1.259 0.493 1.261 0.694 ;
      RECT 1.144 0.493 1.259 0.575 ;
      RECT 1.108 0.255 1.198 0.336 ;
      RECT 1.083 0.693 1.147 0.829 ;
      RECT 1.083 0.281 1.108 0.336 ;
      RECT 1.071 0.281 1.083 0.829 ;
      RECT 1.022 0.281 1.071 0.789 ;
      RECT 0.960 0.175 0.994 0.230 ;
      RECT 0.899 0.175 0.960 0.938 ;
      RECT 0.880 0.657 0.899 0.742 ;
      RECT 0.610 0.811 0.825 0.865 ;
      RECT 0.793 0.338 0.822 0.419 ;
      RECT 0.732 0.338 0.793 0.725 ;
      RECT 0.675 0.670 0.732 0.725 ;
      RECT 0.561 0.939 0.622 1.048 ;
      RECT 0.549 0.368 0.610 0.865 ;
      RECT 0.138 0.939 0.561 0.994 ;
      RECT 0.435 0.368 0.549 0.423 ;
      RECT 0.272 0.699 0.549 0.754 ;
      RECT 0.374 0.336 0.435 0.423 ;
      RECT 0.353 0.161 0.392 0.215 ;
      RECT 0.292 0.161 0.353 0.261 ;
      RECT 0.109 0.206 0.292 0.261 ;
      RECT 0.211 0.657 0.272 0.754 ;
      RECT 0.109 0.874 0.138 0.994 ;
      RECT 0.048 0.206 0.109 0.994 ;
  END
END SEDFFTRX2

MACRO SEDFFHQX2
  CLASS CORE ;
  FOREIGN SEDFFHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.371 0.167 0.511 0.262 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.170 0.490 0.291 0.633 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.862 0.346 5.863 0.733 ;
      RECT 5.803 0.346 5.862 0.767 ;
      RECT 5.758 0.346 5.803 0.427 ;
      RECT 5.763 0.652 5.803 0.767 ;
      RECT 5.758 0.652 5.763 0.733 ;
     END
  END Q

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.772 0.549 1.872 0.693 ;
      RECT 1.702 0.555 1.772 0.610 ;
     END
  END E

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.078 0.433 1.179 0.564 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.448 0.421 2.628 0.512 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.669 -0.080 5.900 0.080 ;
      RECT 5.579 -0.080 5.669 0.122 ;
      RECT 5.294 -0.080 5.579 0.080 ;
      RECT 5.205 -0.080 5.294 0.122 ;
      RECT 4.400 -0.080 5.205 0.080 ;
      RECT 4.311 -0.080 4.400 0.395 ;
      RECT 4.021 -0.080 4.311 0.080 ;
      RECT 3.932 -0.080 4.021 0.342 ;
      RECT 3.430 -0.080 3.932 0.080 ;
      RECT 3.340 -0.080 3.430 0.287 ;
      RECT 2.730 -0.080 3.340 0.080 ;
      RECT 2.641 -0.080 2.730 0.122 ;
      RECT 1.821 -0.080 2.641 0.080 ;
      RECT 1.731 -0.080 1.821 0.122 ;
      RECT 1.113 -0.080 1.731 0.080 ;
      RECT 1.024 -0.080 1.113 0.122 ;
      RECT 0.294 -0.080 1.024 0.080 ;
      RECT 0.205 -0.080 0.294 0.122 ;
      RECT 0.000 -0.080 0.205 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.669 1.120 5.900 1.280 ;
      RECT 5.579 1.078 5.669 1.280 ;
      RECT 5.276 1.120 5.579 1.280 ;
      RECT 5.186 1.078 5.276 1.280 ;
      RECT 3.238 1.120 5.186 1.280 ;
      RECT 3.149 1.078 3.238 1.280 ;
      RECT 2.684 1.120 3.149 1.280 ;
      RECT 2.624 0.902 2.684 1.280 ;
      RECT 1.817 1.120 2.624 1.280 ;
      RECT 1.727 1.078 1.817 1.280 ;
      RECT 1.111 1.120 1.727 1.280 ;
      RECT 1.021 1.078 1.111 1.280 ;
      RECT 0.310 1.120 1.021 1.280 ;
      RECT 0.221 1.078 0.310 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.652 0.500 5.741 0.581 ;
      RECT 5.494 0.526 5.652 0.581 ;
      RECT 5.492 0.292 5.494 0.373 ;
      RECT 5.492 0.526 5.494 0.940 ;
      RECT 5.432 0.292 5.492 0.940 ;
      RECT 5.404 0.292 5.432 0.373 ;
      RECT 5.404 0.748 5.432 0.940 ;
      RECT 5.177 0.855 5.404 0.910 ;
      RECT 5.353 0.543 5.368 0.624 ;
      RECT 5.278 0.543 5.353 0.627 ;
      RECT 5.165 0.573 5.278 0.627 ;
      RECT 5.116 0.683 5.177 0.910 ;
      RECT 5.105 0.213 5.165 0.627 ;
      RECT 5.114 0.855 5.116 0.910 ;
      RECT 5.053 0.855 5.114 1.050 ;
      RECT 5.092 0.213 5.105 0.268 ;
      RECT 5.034 0.573 5.105 0.627 ;
      RECT 5.031 0.174 5.092 0.268 ;
      RECT 3.360 0.995 5.053 1.050 ;
      RECT 4.901 0.330 5.038 0.385 ;
      RECT 4.973 0.573 5.034 0.773 ;
      RECT 4.894 0.174 5.031 0.229 ;
      RECT 4.942 0.718 4.973 0.773 ;
      RECT 4.927 0.718 4.942 0.895 ;
      RECT 4.881 0.718 4.927 0.927 ;
      RECT 4.840 0.330 4.901 0.649 ;
      RECT 4.834 0.150 4.894 0.229 ;
      RECT 4.852 0.814 4.881 0.927 ;
      RECT 4.549 0.873 4.852 0.927 ;
      RECT 4.730 0.594 4.840 0.649 ;
      RECT 4.533 0.150 4.834 0.205 ;
      RECT 4.670 0.737 4.752 0.792 ;
      RECT 4.670 0.261 4.737 0.315 ;
      RECT 4.609 0.261 4.670 0.792 ;
      RECT 4.196 0.470 4.609 0.525 ;
      RECT 4.488 0.735 4.549 0.927 ;
      RECT 4.399 0.594 4.545 0.649 ;
      RECT 4.472 0.150 4.533 0.242 ;
      RECT 4.338 0.594 4.399 0.940 ;
      RECT 3.482 0.886 4.338 0.940 ;
      RECT 4.196 0.276 4.211 0.357 ;
      RECT 4.136 0.276 4.196 0.805 ;
      RECT 4.121 0.276 4.136 0.357 ;
      RECT 4.010 0.508 4.070 0.831 ;
      RECT 3.605 0.776 4.010 0.831 ;
      RECT 3.741 0.289 3.832 0.344 ;
      RECT 3.741 0.665 3.832 0.720 ;
      RECT 3.681 0.289 3.741 0.720 ;
      RECT 3.544 0.231 3.605 0.831 ;
      RECT 3.233 0.554 3.544 0.608 ;
      RECT 3.422 0.843 3.482 0.940 ;
      RECT 3.418 0.357 3.478 0.462 ;
      RECT 2.926 0.843 3.422 0.898 ;
      RECT 3.091 0.357 3.418 0.412 ;
      RECT 3.300 0.954 3.360 1.050 ;
      RECT 2.805 0.954 3.300 1.008 ;
      RECT 3.072 0.268 3.091 0.650 ;
      RECT 3.047 0.255 3.072 0.650 ;
      RECT 3.030 0.255 3.047 0.783 ;
      RECT 2.983 0.255 3.030 0.336 ;
      RECT 2.987 0.595 3.030 0.783 ;
      RECT 2.758 0.394 2.964 0.449 ;
      RECT 2.866 0.665 2.926 0.898 ;
      RECT 2.758 0.665 2.866 0.720 ;
      RECT 2.745 0.776 2.805 1.008 ;
      RECT 2.698 0.257 2.758 0.720 ;
      RECT 2.327 0.776 2.745 0.831 ;
      RECT 2.525 0.257 2.698 0.312 ;
      RECT 2.410 0.665 2.698 0.720 ;
      RECT 2.436 0.231 2.525 0.312 ;
      RECT 1.972 0.982 2.440 1.037 ;
      RECT 2.266 0.306 2.327 0.915 ;
      RECT 2.138 0.390 2.190 0.902 ;
      RECT 2.130 0.306 2.138 0.902 ;
      RECT 2.077 0.306 2.130 0.445 ;
      RECT 2.063 0.833 2.130 0.902 ;
      RECT 2.031 0.542 2.068 0.631 ;
      RECT 1.436 0.833 2.063 0.888 ;
      RECT 2.017 0.150 2.052 0.205 ;
      RECT 2.017 0.542 2.031 0.749 ;
      RECT 1.956 0.150 2.017 0.749 ;
      RECT 1.911 0.954 1.972 1.037 ;
      RECT 1.612 0.192 1.956 0.246 ;
      RECT 1.942 0.668 1.956 0.749 ;
      RECT 0.684 0.954 1.911 1.008 ;
      RECT 1.830 0.375 1.890 0.482 ;
      RECT 1.612 0.427 1.830 0.482 ;
      RECT 1.612 0.668 1.655 0.749 ;
      RECT 1.612 0.302 1.647 0.357 ;
      RECT 1.551 0.161 1.612 0.246 ;
      RECT 1.566 0.302 1.612 0.749 ;
      RECT 1.551 0.302 1.566 0.736 ;
      RECT 1.298 0.161 1.551 0.215 ;
      RECT 1.520 0.526 1.551 0.613 ;
      RECT 1.436 0.287 1.450 0.368 ;
      RECT 1.375 0.287 1.436 0.899 ;
      RECT 1.361 0.287 1.375 0.368 ;
      RECT 1.007 0.844 1.375 0.899 ;
      RECT 1.261 0.300 1.300 0.725 ;
      RECT 1.240 0.287 1.261 0.738 ;
      RECT 1.171 0.287 1.240 0.368 ;
      RECT 1.171 0.657 1.240 0.738 ;
      RECT 0.947 0.202 1.007 0.899 ;
      RECT 0.889 0.202 0.947 0.257 ;
      RECT 0.797 0.844 0.947 0.899 ;
      RECT 0.828 0.163 0.889 0.257 ;
      RECT 0.824 0.318 0.885 0.733 ;
      RECT 0.797 0.163 0.828 0.218 ;
      RECT 0.785 0.469 0.824 0.554 ;
      RECT 0.686 0.343 0.715 0.424 ;
      RECT 0.669 0.343 0.686 0.501 ;
      RECT 0.669 0.820 0.684 1.008 ;
      RECT 0.626 0.343 0.669 1.008 ;
      RECT 0.623 0.446 0.626 1.008 ;
      RECT 0.609 0.446 0.623 0.901 ;
      RECT 0.594 0.820 0.609 0.901 ;
      RECT 0.530 0.969 0.544 1.050 ;
      RECT 0.455 0.935 0.530 1.050 ;
      RECT 0.476 0.343 0.505 0.424 ;
      RECT 0.476 0.746 0.484 0.827 ;
      RECT 0.415 0.343 0.476 0.827 ;
      RECT 0.137 0.935 0.455 0.989 ;
      RECT 0.394 0.746 0.415 0.827 ;
      RECT 0.108 0.343 0.137 0.424 ;
      RECT 0.108 0.746 0.137 0.989 ;
      RECT 0.076 0.343 0.108 0.989 ;
      RECT 0.047 0.343 0.076 0.827 ;
  END
END SEDFFHQX2

MACRO SDFFSX2
  CLASS CORE ;
  FOREIGN SDFFSX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.197 0.951 3.307 1.033 ;
      RECT 2.968 0.951 3.197 1.006 ;
      RECT 2.907 0.951 2.968 1.026 ;
      RECT 2.688 0.971 2.907 1.026 ;
      RECT 2.627 0.954 2.688 1.026 ;
      RECT 1.904 0.954 2.627 1.008 ;
      RECT 1.843 0.954 1.904 1.010 ;
      RECT 1.828 0.955 1.843 1.010 ;
     END
  END SN

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.741 0.475 0.881 0.633 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.213 0.433 0.441 0.500 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.955 0.295 3.991 0.361 ;
      RECT 3.893 0.163 3.955 0.707 ;
      RECT 3.811 0.163 3.893 0.218 ;
      RECT 3.867 0.652 3.893 0.707 ;
      RECT 3.776 0.652 3.867 0.733 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.285 0.315 4.343 0.749 ;
      RECT 4.281 0.177 4.285 0.749 ;
      RECT 4.195 0.177 4.281 0.370 ;
      RECT 4.251 0.694 4.281 0.767 ;
      RECT 4.160 0.694 4.251 0.999 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.112 0.433 1.203 0.595 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.674 0.219 0.767 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.079 -0.080 4.400 0.080 ;
      RECT 4.017 -0.080 4.079 0.224 ;
      RECT 3.565 -0.080 4.017 0.080 ;
      RECT 3.475 -0.080 3.565 0.122 ;
      RECT 3.080 -0.080 3.475 0.080 ;
      RECT 2.989 -0.080 3.080 0.246 ;
      RECT 2.401 -0.080 2.989 0.080 ;
      RECT 2.340 -0.080 2.401 0.328 ;
      RECT 1.808 -0.080 2.340 0.080 ;
      RECT 1.717 -0.080 1.808 0.254 ;
      RECT 0.956 -0.080 1.717 0.080 ;
      RECT 0.865 -0.080 0.956 0.122 ;
      RECT 0.380 -0.080 0.865 0.080 ;
      RECT 0.289 -0.080 0.380 0.122 ;
      RECT 0.000 -0.080 0.289 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.059 1.120 4.400 1.280 ;
      RECT 3.968 0.942 4.059 1.280 ;
      RECT 3.531 1.120 3.968 1.280 ;
      RECT 3.440 0.835 3.531 1.280 ;
      RECT 3.136 1.120 3.440 1.280 ;
      RECT 3.045 1.078 3.136 1.280 ;
      RECT 2.532 1.120 3.045 1.280 ;
      RECT 2.384 1.078 2.532 1.280 ;
      RECT 2.139 1.120 2.384 1.280 ;
      RECT 2.048 1.078 2.139 1.280 ;
      RECT 1.765 1.120 2.048 1.280 ;
      RECT 1.675 1.078 1.765 1.280 ;
      RECT 0.944 1.120 1.675 1.280 ;
      RECT 0.853 0.957 0.944 1.280 ;
      RECT 0.288 1.120 0.853 1.280 ;
      RECT 0.197 1.078 0.288 1.280 ;
      RECT 0.000 1.120 0.197 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.099 0.493 4.157 0.574 ;
      RECT 4.037 0.493 4.099 0.844 ;
      RECT 3.723 0.789 4.037 0.844 ;
      RECT 3.715 0.320 3.757 0.401 ;
      RECT 3.715 0.789 3.723 0.901 ;
      RECT 3.653 0.320 3.715 0.901 ;
      RECT 3.632 0.820 3.653 0.901 ;
      RECT 3.553 0.480 3.583 0.561 ;
      RECT 3.492 0.315 3.553 0.755 ;
      RECT 3.421 0.315 3.492 0.370 ;
      RECT 3.339 0.700 3.492 0.755 ;
      RECT 3.331 0.300 3.421 0.381 ;
      RECT 3.375 0.521 3.403 0.602 ;
      RECT 3.312 0.521 3.375 0.636 ;
      RECT 3.248 0.700 3.339 0.893 ;
      RECT 2.999 0.315 3.331 0.370 ;
      RECT 2.812 0.581 3.312 0.636 ;
      RECT 2.937 0.315 2.999 0.525 ;
      RECT 2.908 0.444 2.937 0.525 ;
      RECT 2.812 0.324 2.813 0.405 ;
      RECT 2.751 0.324 2.812 0.917 ;
      RECT 2.723 0.324 2.751 0.405 ;
      RECT 2.623 0.605 2.684 0.899 ;
      RECT 2.547 0.445 2.661 0.526 ;
      RECT 1.665 0.844 2.623 0.899 ;
      RECT 2.485 0.398 2.547 0.719 ;
      RECT 2.279 0.398 2.485 0.452 ;
      RECT 2.341 0.664 2.485 0.719 ;
      RECT 2.156 0.510 2.424 0.590 ;
      RECT 2.251 0.664 2.341 0.745 ;
      RECT 2.217 0.173 2.279 0.452 ;
      RECT 2.008 0.173 2.217 0.227 ;
      RECT 2.095 0.343 2.156 0.769 ;
      RECT 1.723 0.714 2.095 0.769 ;
      RECT 1.848 0.582 2.019 0.637 ;
      RECT 1.917 0.151 2.008 0.227 ;
      RECT 1.787 0.463 1.848 0.637 ;
      RECT 1.517 0.463 1.787 0.518 ;
      RECT 1.661 0.575 1.723 0.769 ;
      RECT 1.604 0.844 1.665 0.973 ;
      RECT 1.632 0.575 1.661 0.656 ;
      RECT 1.460 0.918 1.604 0.973 ;
      RECT 1.517 0.181 1.532 0.262 ;
      RECT 1.456 0.181 1.517 0.782 ;
      RECT 1.399 0.918 1.460 1.049 ;
      RECT 1.441 0.181 1.456 0.262 ;
      RECT 1.391 0.701 1.456 0.782 ;
      RECT 1.329 0.994 1.399 1.049 ;
      RECT 1.329 0.358 1.379 0.465 ;
      RECT 1.268 0.358 1.329 1.049 ;
      RECT 1.228 0.181 1.319 0.262 ;
      RECT 1.067 0.994 1.268 1.049 ;
      RECT 0.704 0.194 1.228 0.249 ;
      RECT 1.132 0.723 1.193 0.939 ;
      RECT 0.647 0.723 1.132 0.777 ;
      RECT 1.005 0.832 1.067 1.049 ;
      RECT 0.940 0.308 1.031 0.389 ;
      RECT 0.792 0.832 1.005 0.887 ;
      RECT 0.659 0.321 0.940 0.376 ;
      RECT 0.731 0.832 0.792 1.039 ;
      RECT 0.449 0.985 0.731 1.039 ;
      RECT 0.643 0.165 0.704 0.249 ;
      RECT 0.597 0.321 0.659 0.656 ;
      RECT 0.585 0.723 0.647 0.929 ;
      RECT 0.503 0.165 0.643 0.220 ;
      RECT 0.503 0.321 0.597 0.402 ;
      RECT 0.568 0.575 0.597 0.656 ;
      RECT 0.544 0.848 0.585 0.929 ;
      RECT 0.501 0.601 0.568 0.656 ;
      RECT 0.440 0.601 0.501 0.752 ;
      RECT 0.388 0.856 0.449 1.039 ;
      RECT 0.411 0.671 0.440 0.752 ;
      RECT 0.341 0.856 0.388 0.911 ;
      RECT 0.280 0.560 0.341 0.911 ;
      RECT 0.109 0.560 0.280 0.614 ;
      RECT 0.139 0.843 0.280 0.911 ;
      RECT 0.109 0.293 0.139 0.374 ;
      RECT 0.048 0.830 0.139 0.911 ;
      RECT 0.048 0.293 0.109 0.614 ;
  END
END SDFFSX2

MACRO SDFFRHQX2
  CLASS CORE ;
  FOREIGN SDFFRHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.865 0.567 0.984 0.629 ;
      RECT 0.776 0.548 0.865 0.629 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.383 0.415 0.491 0.543 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.216 0.632 4.357 0.763 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.937 0.275 4.998 0.729 ;
      RECT 4.643 0.275 4.937 0.330 ;
      RECT 4.817 0.674 4.937 0.729 ;
      RECT 4.727 0.674 4.817 0.960 ;
      RECT 4.641 0.225 4.643 0.330 ;
      RECT 4.551 0.151 4.641 0.344 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.019 0.418 1.177 0.510 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.290 0.506 0.310 0.617 ;
      RECT 0.230 0.506 0.290 0.627 ;
      RECT 0.158 0.506 0.230 0.617 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.840 -0.080 5.200 0.080 ;
      RECT 4.751 -0.080 4.840 0.122 ;
      RECT 4.382 -0.080 4.751 0.080 ;
      RECT 4.135 -0.080 4.382 0.122 ;
      RECT 3.782 -0.080 4.135 0.080 ;
      RECT 3.693 -0.080 3.782 0.122 ;
      RECT 2.754 -0.080 3.693 0.080 ;
      RECT 2.664 -0.080 2.754 0.292 ;
      RECT 1.731 -0.080 2.664 0.080 ;
#      RECT 2.035 0.303 2.125 0.359 ;
#      RECT 1.731 0.303 2.035 0.353 ;
      RECT 1.670 -0.080 1.731 0.328 ;
      RECT 1.641 -0.080 1.670 0.327 ;
      RECT 0.826 -0.080 1.641 0.080 ;
      RECT 0.737 -0.080 0.826 0.122 ;
      RECT 0.284 -0.080 0.737 0.080 ;
      RECT 0.194 -0.080 0.284 0.122 ;
      RECT 0.000 -0.080 0.194 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.153 1.120 5.200 1.280 ;
      RECT 5.063 0.800 5.153 1.280 ;
      RECT 4.457 1.120 5.063 1.280 ;
      RECT 4.367 1.078 4.457 1.280 ;
      RECT 4.089 1.120 4.367 1.280 ;
      RECT 4.000 1.078 4.089 1.280 ;
      RECT 3.778 1.120 4.000 1.280 ;
      RECT 3.662 1.078 3.778 1.280 ;
      RECT 2.759 1.120 3.662 1.280 ;
      RECT 2.670 1.078 2.759 1.280 ;
      RECT 1.754 1.120 2.670 1.280 ;
      RECT 1.665 0.997 1.754 1.280 ;
      RECT 0.919 1.120 1.665 1.280 ;
      RECT 0.830 1.001 0.919 1.280 ;
      RECT 0.347 1.120 0.830 1.280 ;
      RECT 0.336 1.013 0.347 1.280 ;
      RECT 0.247 0.972 0.336 1.280 ;
      RECT 0.236 1.013 0.247 1.280 ;
      RECT 0.000 1.120 0.236 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.725 0.538 4.877 0.619 ;
      RECT 4.664 0.399 4.725 0.619 ;
      RECT 4.411 0.399 4.664 0.454 ;
      RECT 4.473 0.523 4.562 0.612 ;
      RECT 4.289 0.523 4.473 0.577 ;
      RECT 4.350 0.206 4.411 0.454 ;
      RECT 3.925 0.206 4.350 0.261 ;
      RECT 4.226 0.838 4.315 0.919 ;
      RECT 4.199 0.352 4.289 0.577 ;
      RECT 4.025 0.838 4.226 0.893 ;
      RECT 4.094 0.523 4.199 0.577 ;
      RECT 4.025 0.517 4.094 0.598 ;
      RECT 4.005 0.517 4.025 0.994 ;
      RECT 3.921 0.336 4.010 0.417 ;
      RECT 3.964 0.543 4.005 0.994 ;
      RECT 3.431 0.939 3.964 0.994 ;
      RECT 3.832 0.206 3.925 0.273 ;
      RECT 3.807 0.349 3.921 0.404 ;
      RECT 3.425 0.206 3.832 0.261 ;
      RECT 3.807 0.736 3.821 0.817 ;
      RECT 3.746 0.349 3.807 0.817 ;
      RECT 3.732 0.605 3.746 0.817 ;
      RECT 3.658 0.605 3.732 0.686 ;
      RECT 3.484 0.360 3.498 0.440 ;
      RECT 3.459 0.360 3.484 0.688 ;
      RECT 3.423 0.360 3.459 0.714 ;
      RECT 3.371 0.939 3.431 1.039 ;
      RECT 3.334 0.170 3.425 0.261 ;
      RECT 3.409 0.360 3.423 0.440 ;
      RECT 3.369 0.633 3.423 0.714 ;
      RECT 2.916 0.985 3.371 1.039 ;
      RECT 3.310 0.795 3.362 0.876 ;
      RECT 3.158 0.206 3.334 0.261 ;
      RECT 3.305 0.338 3.325 0.419 ;
      RECT 3.305 0.795 3.310 0.915 ;
      RECT 3.245 0.338 3.305 0.915 ;
      RECT 3.236 0.338 3.245 0.419 ;
      RECT 3.037 0.861 3.245 0.915 ;
      RECT 3.098 0.206 3.158 0.786 ;
      RECT 3.058 0.206 3.098 0.419 ;
      RECT 2.983 0.817 3.037 0.915 ;
      RECT 2.977 0.804 2.983 0.915 ;
      RECT 2.968 0.804 2.977 0.885 ;
      RECT 2.943 0.362 2.968 0.885 ;
      RECT 2.907 0.240 2.943 0.885 ;
      RECT 2.856 0.939 2.916 1.039 ;
      RECT 2.853 0.240 2.907 0.417 ;
      RECT 2.894 0.804 2.907 0.885 ;
      RECT 2.621 0.817 2.894 0.871 ;
      RECT 2.184 0.939 2.856 0.994 ;
      RECT 2.550 0.362 2.853 0.417 ;
      RECT 2.786 0.471 2.847 0.746 ;
      RECT 2.428 0.471 2.786 0.526 ;
      RECT 2.437 0.692 2.786 0.746 ;
      RECT 2.307 0.582 2.684 0.637 ;
      RECT 2.532 0.802 2.621 0.883 ;
      RECT 2.490 0.252 2.550 0.417 ;
      RECT 2.377 0.692 2.437 0.829 ;
      RECT 2.368 0.319 2.428 0.526 ;
      RECT 2.348 0.748 2.377 0.829 ;
      RECT 2.336 0.319 2.368 0.374 ;
      RECT 2.307 0.293 2.336 0.374 ;
      RECT 2.247 0.176 2.307 0.374 ;
      RECT 2.247 0.477 2.307 0.637 ;
      RECT 1.901 0.176 2.247 0.231 ;
      RECT 1.976 0.477 2.247 0.532 ;
      RECT 2.123 0.607 2.184 0.994 ;
      RECT 1.916 0.477 1.976 0.876 ;
      RECT 1.915 0.477 1.916 0.532 ;
      RECT 1.853 0.795 1.916 0.876 ;
      RECT 1.825 0.398 1.915 0.532 ;
      RECT 1.812 0.150 1.901 0.231 ;
      RECT 1.743 0.607 1.832 0.701 ;
      RECT 1.656 0.477 1.825 0.532 ;
      RECT 1.454 0.646 1.743 0.701 ;
      RECT 1.595 0.477 1.656 0.590 ;
      RECT 1.567 0.510 1.595 0.590 ;
      RECT 1.494 0.902 1.509 0.983 ;
      RECT 1.419 0.901 1.494 0.983 ;
      RECT 1.393 0.176 1.454 0.792 ;
      RECT 1.299 0.901 1.419 0.956 ;
      RECT 1.372 0.176 1.393 0.231 ;
      RECT 1.359 0.698 1.393 0.792 ;
      RECT 1.283 0.150 1.372 0.231 ;
      RECT 1.299 0.445 1.301 0.630 ;
      RECT 1.241 0.445 1.299 0.956 ;
      RECT 1.238 0.575 1.241 0.956 ;
      RECT 0.599 0.732 1.238 0.787 ;
      RECT 1.098 0.202 1.187 0.283 ;
      RECT 1.117 0.856 1.178 0.995 ;
      RECT 0.755 0.856 1.117 0.911 ;
      RECT 0.545 0.206 1.098 0.261 ;
      RECT 0.852 0.324 0.901 0.405 ;
      RECT 0.624 0.323 0.852 0.405 ;
      RECT 0.695 0.856 0.755 0.993 ;
      RECT 0.615 0.938 0.695 0.993 ;
      RECT 0.624 0.595 0.688 0.676 ;
      RECT 0.599 0.323 0.624 0.676 ;
      RECT 0.525 0.938 0.615 1.019 ;
      RECT 0.552 0.323 0.599 0.663 ;
      RECT 0.538 0.732 0.599 0.858 ;
      RECT 0.469 0.608 0.552 0.663 ;
      RECT 0.485 0.165 0.545 0.261 ;
      RECT 0.137 0.804 0.538 0.858 ;
      RECT 0.378 0.165 0.485 0.220 ;
      RECT 0.408 0.608 0.469 0.748 ;
      RECT 0.122 0.318 0.137 0.399 ;
      RECT 0.097 0.671 0.137 0.864 ;
      RECT 0.097 0.318 0.122 0.450 ;
      RECT 0.047 0.318 0.097 0.864 ;
      RECT 0.037 0.395 0.047 0.726 ;
  END
END SDFFRHQX2

MACRO SDFFRX2
  CLASS CORE ;
  FOREIGN SDFFRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.743 0.538 0.902 0.638 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.450 0.295 0.471 0.371 ;
      RECT 0.450 0.460 0.465 0.540 ;
      RECT 0.390 0.295 0.450 0.540 ;
      RECT 0.376 0.460 0.390 0.540 ;
     END
  END SE

  PIN RN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.903 0.685 1.917 0.807 ;
      RECT 1.828 0.656 1.903 0.807 ;
      RECT 1.790 0.656 1.828 0.794 ;
      RECT 1.778 0.685 1.790 0.771 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.781 0.435 4.797 0.494 ;
      RECT 4.781 0.698 4.796 0.779 ;
      RECT 4.733 0.435 4.781 0.779 ;
      RECT 4.721 0.326 4.733 0.779 ;
      RECT 4.672 0.326 4.721 0.489 ;
      RECT 4.706 0.698 4.721 0.779 ;
      RECT 4.643 0.326 4.672 0.407 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.142 0.227 5.159 0.769 ;
      RECT 5.140 0.227 5.142 0.779 ;
      RECT 5.081 0.163 5.140 0.779 ;
      RECT 5.050 0.163 5.081 0.387 ;
      RECT 5.053 0.693 5.081 0.779 ;
      RECT 5.045 0.698 5.053 0.779 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.008 0.369 1.177 0.505 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.253 0.429 0.302 0.505 ;
      RECT 0.164 0.408 0.253 0.671 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.920 -0.080 5.200 0.080 ;
      RECT 4.860 -0.080 4.920 0.355 ;
      RECT 4.402 -0.080 4.860 0.080 ;
      RECT 4.312 -0.080 4.402 0.268 ;
      RECT 4.010 -0.080 4.312 0.080 ;
      RECT 3.921 -0.080 4.010 0.122 ;
      RECT 3.522 -0.080 3.921 0.080 ;
      RECT 3.433 -0.080 3.522 0.283 ;
      RECT 2.805 -0.080 3.433 0.080 ;
      RECT 2.716 -0.080 2.805 0.311 ;
      RECT 2.358 -0.080 2.716 0.080 ;
      RECT 2.269 -0.080 2.358 0.214 ;
      RECT 2.038 -0.080 2.269 0.090 ;
      RECT 1.926 -0.080 2.038 0.303 ;
      RECT 0.825 -0.080 1.926 0.080 ;
      RECT 0.735 -0.080 0.825 0.122 ;
      RECT 0.284 -0.080 0.735 0.080 ;
      RECT 0.194 -0.080 0.284 0.122 ;
      RECT 0.000 -0.080 0.194 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.964 1.120 5.200 1.280 ;
      RECT 4.874 0.986 4.964 1.280 ;
      RECT 4.423 1.120 4.874 1.280 ;
      RECT 4.333 0.891 4.423 1.280 ;
      RECT 3.693 1.120 4.333 1.280 ;
      RECT 3.603 0.986 3.693 1.280 ;
      RECT 2.979 1.120 3.603 1.280 ;
      RECT 2.600 1.047 2.979 1.280 ;
      RECT 1.838 1.120 2.600 1.280 ;
      RECT 1.749 1.078 1.838 1.280 ;
      RECT 1.008 1.120 1.749 1.280 ;
      RECT 0.919 0.963 1.008 1.280 ;
      RECT 0.284 1.120 0.919 1.280 ;
      RECT 0.194 1.078 0.284 1.280 ;
      RECT 0.000 1.120 0.194 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.960 0.455 5.020 0.632 ;
      RECT 4.948 0.577 4.960 0.632 ;
      RECT 4.887 0.577 4.948 0.906 ;
      RECT 4.612 0.851 4.887 0.906 ;
      RECT 4.583 0.851 4.612 0.957 ;
      RECT 4.583 0.158 4.601 0.239 ;
      RECT 4.522 0.158 4.583 0.957 ;
      RECT 4.512 0.158 4.522 0.239 ;
      RECT 4.448 0.379 4.462 0.487 ;
      RECT 4.387 0.379 4.448 0.754 ;
      RECT 4.373 0.379 4.387 0.487 ;
      RECT 4.244 0.699 4.387 0.754 ;
      RECT 4.213 0.432 4.373 0.487 ;
      RECT 4.184 0.699 4.244 0.836 ;
      RECT 4.152 0.217 4.213 0.487 ;
      RECT 4.039 0.781 4.184 0.836 ;
      RECT 4.123 0.217 4.152 0.298 ;
      RECT 3.974 0.432 4.152 0.487 ;
      RECT 4.010 0.781 4.039 0.862 ;
      RECT 3.950 0.781 4.010 1.017 ;
      RECT 3.858 0.586 3.989 0.667 ;
      RECT 3.899 0.388 3.974 0.487 ;
      RECT 3.876 0.936 3.950 1.017 ;
      RECT 3.884 0.388 3.899 0.469 ;
      RECT 3.824 0.586 3.858 0.794 ;
      RECT 3.763 0.401 3.824 0.794 ;
      RECT 3.737 0.401 3.763 0.456 ;
      RECT 3.761 0.638 3.763 0.794 ;
      RECT 3.494 0.739 3.761 0.794 ;
      RECT 3.677 0.292 3.737 0.456 ;
      RECT 3.689 0.525 3.703 0.580 ;
      RECT 3.628 0.525 3.689 0.581 ;
      RECT 3.616 0.292 3.677 0.418 ;
      RECT 3.526 0.526 3.628 0.581 ;
      RECT 3.178 0.363 3.616 0.418 ;
      RECT 3.465 0.473 3.526 0.581 ;
      RECT 3.434 0.739 3.494 0.829 ;
      RECT 3.057 0.473 3.465 0.527 ;
      RECT 3.346 0.774 3.434 0.829 ;
      RECT 3.257 0.774 3.346 0.855 ;
      RECT 3.194 0.619 3.283 0.700 ;
      RECT 3.190 0.645 3.194 0.700 ;
      RECT 3.129 0.645 3.190 0.929 ;
      RECT 3.117 0.260 3.178 0.418 ;
      RECT 2.630 0.874 3.129 0.929 ;
      RECT 3.073 0.260 3.117 0.340 ;
      RECT 2.997 0.406 3.057 0.818 ;
      RECT 2.595 0.406 2.997 0.461 ;
      RECT 2.750 0.763 2.997 0.818 ;
      RECT 2.847 0.517 2.936 0.687 ;
      RECT 2.420 0.517 2.847 0.571 ;
      RECT 2.671 0.626 2.760 0.707 ;
      RECT 2.630 0.639 2.671 0.707 ;
      RECT 2.570 0.639 2.630 0.929 ;
      RECT 2.593 0.287 2.595 0.461 ;
      RECT 2.565 0.274 2.593 0.461 ;
      RECT 2.515 0.874 2.570 0.929 ;
      RECT 2.519 0.158 2.565 0.461 ;
      RECT 2.504 0.158 2.519 0.355 ;
      RECT 2.454 0.874 2.515 1.037 ;
      RECT 2.435 0.158 2.504 0.213 ;
      RECT 1.961 0.982 2.454 1.037 ;
      RECT 2.360 0.375 2.420 0.758 ;
      RECT 2.227 0.375 2.360 0.430 ;
      RECT 2.310 0.704 2.360 0.758 ;
      RECT 2.310 0.826 2.324 0.907 ;
      RECT 2.249 0.704 2.310 0.907 ;
      RECT 2.210 0.510 2.299 0.590 ;
      RECT 2.235 0.826 2.249 0.907 ;
      RECT 2.167 0.346 2.227 0.430 ;
      RECT 2.097 0.523 2.210 0.577 ;
      RECT 2.138 0.346 2.167 0.427 ;
      RECT 1.660 0.373 2.138 0.427 ;
      RECT 2.097 0.845 2.112 0.926 ;
      RECT 2.037 0.523 2.097 0.926 ;
      RECT 2.035 0.523 2.037 0.577 ;
      RECT 2.022 0.845 2.037 0.926 ;
      RECT 1.891 0.483 2.035 0.577 ;
      RECT 1.900 0.939 1.961 1.037 ;
      RECT 1.666 0.939 1.900 0.994 ;
      RECT 1.765 0.161 1.854 0.264 ;
      RECT 1.488 0.161 1.765 0.215 ;
      RECT 1.606 0.939 1.666 1.013 ;
      RECT 1.573 0.373 1.660 0.496 ;
      RECT 1.366 0.958 1.606 1.013 ;
      RECT 1.571 0.415 1.573 0.496 ;
      RECT 1.493 0.786 1.507 0.867 ;
      RECT 1.488 0.781 1.493 0.867 ;
      RECT 1.427 0.161 1.488 0.867 ;
      RECT 1.303 0.221 1.427 0.302 ;
      RECT 1.418 0.786 1.427 0.867 ;
      RECT 1.339 0.945 1.366 1.026 ;
      RECT 1.328 0.394 1.339 1.026 ;
      RECT 1.279 0.381 1.328 1.026 ;
      RECT 1.238 0.381 1.279 0.462 ;
      RECT 1.276 0.945 1.279 1.026 ;
      RECT 1.152 0.945 1.276 1.000 ;
      RECT 1.104 0.679 1.194 0.760 ;
      RECT 1.093 0.206 1.182 0.302 ;
      RECT 1.091 0.821 1.152 1.000 ;
      RECT 0.650 0.699 1.104 0.754 ;
      RECT 0.674 0.206 1.093 0.261 ;
      RECT 0.661 0.821 1.091 0.876 ;
      RECT 0.793 0.389 0.882 0.470 ;
      RECT 0.633 0.402 0.793 0.457 ;
      RECT 0.613 0.158 0.674 0.261 ;
      RECT 0.600 0.821 0.661 1.008 ;
      RECT 0.586 0.348 0.633 0.493 ;
      RECT 0.469 0.158 0.613 0.213 ;
      RECT 0.137 0.954 0.600 1.008 ;
      RECT 0.544 0.348 0.586 0.652 ;
      RECT 0.542 0.438 0.544 0.652 ;
      RECT 0.525 0.438 0.542 0.757 ;
      RECT 0.494 0.596 0.525 0.757 ;
      RECT 0.482 0.596 0.494 0.898 ;
      RECT 0.433 0.676 0.482 0.898 ;
      RECT 0.378 0.158 0.469 0.229 ;
      RECT 0.404 0.817 0.433 0.898 ;
      RECT 0.104 0.262 0.137 0.343 ;
      RECT 0.104 0.864 0.137 1.008 ;
      RECT 0.043 0.262 0.104 1.008 ;
  END
END SDFFRX2

MACRO SDFFHQX2
  CLASS CORE ;
  FOREIGN SDFFHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.790 0.433 0.838 0.500 ;
      RECT 0.655 0.412 0.790 0.500 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.059 0.648 1.088 0.729 ;
      RECT 0.998 0.574 1.059 0.729 ;
      RECT 0.663 0.574 0.998 0.629 ;
      RECT 0.562 0.567 0.663 0.635 ;
      RECT 0.544 0.568 0.562 0.635 ;
     END
  END SE

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.855 0.167 3.945 0.248 ;
      RECT 3.756 0.193 3.855 0.248 ;
      RECT 3.756 0.700 3.813 0.767 ;
      RECT 3.695 0.193 3.756 0.767 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.051 0.335 1.184 0.494 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.512 0.327 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.147 -0.080 4.200 0.080 ;
      RECT 4.057 -0.080 4.147 0.211 ;
      RECT 3.733 -0.080 4.057 0.080 ;
      RECT 3.643 -0.080 3.733 0.122 ;
      RECT 3.199 -0.080 3.643 0.080 ;
      RECT 3.138 -0.080 3.199 0.241 ;
      RECT 2.376 -0.080 3.138 0.080 ;
      RECT 2.286 -0.080 2.376 0.308 ;
      RECT 1.766 -0.080 2.286 0.080 ;
      RECT 1.676 -0.080 1.766 0.287 ;
      RECT 0.833 -0.080 1.676 0.080 ;
      RECT 0.742 -0.080 0.833 0.122 ;
      RECT 0.321 -0.080 0.742 0.080 ;
      RECT 0.321 0.358 0.329 0.409 ;
      RECT 0.231 -0.080 0.321 0.409 ;
      RECT 0.000 -0.080 0.231 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.972 1.120 4.200 1.280 ;
      RECT 3.882 1.078 3.972 1.280 ;
      RECT 3.447 1.120 3.882 1.280 ;
      RECT 2.983 1.078 3.447 1.280 ;
      RECT 2.272 1.120 2.983 1.280 ;
      RECT 2.182 1.078 2.272 1.280 ;
      RECT 1.087 1.120 2.182 1.280 ;
      RECT 0.997 1.065 1.087 1.280 ;
      RECT 0.403 1.120 0.997 1.280 ;
      RECT 0.313 1.078 0.403 1.280 ;
      RECT 0.000 1.120 0.313 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.997 0.374 4.058 0.986 ;
      RECT 3.945 0.374 3.997 0.429 ;
      RECT 3.770 0.931 3.997 0.986 ;
      RECT 3.855 0.348 3.945 0.429 ;
      RECT 3.874 0.544 3.935 0.876 ;
      RECT 3.634 0.821 3.874 0.876 ;
      RECT 3.679 0.931 3.770 1.040 ;
      RECT 3.458 0.931 3.679 0.986 ;
      RECT 3.573 0.357 3.634 0.876 ;
      RECT 3.426 0.357 3.573 0.412 ;
      RECT 3.206 0.800 3.573 0.855 ;
      RECT 3.451 0.467 3.512 0.745 ;
      RECT 3.367 0.917 3.458 0.998 ;
      RECT 2.945 0.467 3.451 0.521 ;
      RECT 2.872 0.690 3.451 0.745 ;
      RECT 3.336 0.277 3.426 0.412 ;
      RECT 2.681 0.576 3.370 0.631 ;
      RECT 3.066 0.357 3.336 0.412 ;
      RECT 3.177 0.800 3.206 0.881 ;
      RECT 3.116 0.800 3.177 0.998 ;
      RECT 2.681 0.943 3.116 0.998 ;
      RECT 3.005 0.152 3.066 0.412 ;
      RECT 2.770 0.152 3.005 0.207 ;
      RECT 2.884 0.262 2.945 0.521 ;
      RECT 2.577 0.344 2.884 0.399 ;
      RECT 2.811 0.690 2.872 0.888 ;
      RECT 2.781 0.807 2.811 0.888 ;
      RECT 2.475 0.807 2.781 0.862 ;
      RECT 2.709 0.152 2.770 0.289 ;
      RECT 2.678 0.235 2.709 0.289 ;
      RECT 2.652 0.576 2.681 0.752 ;
      RECT 2.591 0.917 2.681 0.998 ;
      RECT 2.591 0.454 2.652 0.752 ;
      RECT 2.161 0.454 2.591 0.508 ;
      RECT 2.353 0.698 2.591 0.752 ;
      RECT 2.516 0.262 2.577 0.399 ;
      RECT 2.487 0.262 2.516 0.343 ;
      RECT 2.414 0.807 2.475 0.888 ;
      RECT 2.231 0.563 2.453 0.618 ;
      RECT 2.292 0.698 2.353 1.008 ;
      RECT 1.678 0.954 2.292 1.008 ;
      RECT 2.170 0.563 2.231 0.899 ;
      RECT 1.963 0.844 2.170 0.899 ;
      RECT 2.125 0.263 2.164 0.344 ;
      RECT 2.100 0.150 2.125 0.344 ;
      RECT 2.100 0.563 2.109 0.706 ;
      RECT 2.048 0.150 2.100 0.706 ;
      RECT 2.039 0.150 2.048 0.618 ;
      RECT 2.030 0.150 2.039 0.205 ;
      RECT 1.902 0.226 1.963 0.899 ;
      RECT 1.661 0.514 1.902 0.595 ;
      RECT 1.600 0.368 1.808 0.423 ;
      RECT 1.677 0.933 1.678 1.019 ;
      RECT 1.588 0.926 1.677 1.019 ;
      RECT 1.539 0.368 1.600 0.857 ;
      RECT 1.478 0.926 1.588 0.988 ;
      RECT 1.488 0.368 1.539 0.423 ;
      RECT 1.427 0.219 1.488 0.423 ;
      RECT 1.417 0.619 1.478 0.988 ;
      RECT 1.405 0.219 1.427 0.274 ;
      RECT 1.343 0.619 1.417 0.674 ;
      RECT 0.936 0.933 1.417 0.988 ;
      RECT 1.315 0.193 1.405 0.274 ;
      RECT 1.266 0.769 1.356 0.850 ;
      RECT 1.343 0.329 1.344 0.410 ;
      RECT 1.282 0.329 1.343 0.674 ;
      RECT 1.254 0.329 1.282 0.410 ;
      RECT 0.814 0.795 1.266 0.850 ;
      RECT 1.103 0.179 1.193 0.260 ;
      RECT 0.677 0.193 1.103 0.248 ;
      RECT 0.851 0.302 0.941 0.373 ;
      RECT 0.875 0.933 0.936 1.050 ;
      RECT 0.525 0.995 0.875 1.050 ;
      RECT 0.562 0.302 0.851 0.357 ;
      RECT 0.753 0.795 0.814 0.936 ;
      RECT 0.609 0.881 0.753 0.936 ;
      RECT 0.602 0.724 0.692 0.805 ;
      RECT 0.616 0.154 0.677 0.248 ;
      RECT 0.382 0.154 0.616 0.208 ;
      RECT 0.552 0.724 0.602 0.779 ;
      RECT 0.487 0.302 0.562 0.424 ;
      RECT 0.451 0.700 0.552 0.779 ;
      RECT 0.464 0.858 0.525 1.050 ;
      RECT 0.472 0.343 0.487 0.424 ;
      RECT 0.451 0.369 0.472 0.424 ;
      RECT 0.209 0.858 0.464 0.913 ;
      RECT 0.419 0.369 0.451 0.779 ;
      RECT 0.390 0.369 0.419 0.755 ;
      RECT 0.151 0.719 0.209 0.913 ;
      RECT 0.103 0.319 0.151 0.913 ;
      RECT 0.090 0.319 0.103 0.788 ;
      RECT 0.048 0.319 0.090 0.400 ;

      LAYER Metal2 ;
      RECT 0.200 0.225 2.340 0.275 ;
      RECT 2.500 0.525 4.000 0.575 ;
      RECT 0.200 0.825 3.040 0.875 ;
  END
END SDFFHQX2

MACRO SDFFX2
  CLASS CORE ;
  FOREIGN SDFFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN SI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.765 0.433 0.843 0.500 ;
      RECT 0.672 0.412 0.765 0.500 ;
     END
  END SI

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.081 0.648 1.111 0.729 ;
      RECT 1.020 0.573 1.081 0.729 ;
      RECT 1.019 0.573 1.020 0.633 ;
      RECT 0.667 0.573 1.019 0.627 ;
      RECT 0.547 0.567 0.667 0.633 ;
     END
  END SE

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.105 0.323 4.167 0.793 ;
      RECT 4.085 0.323 4.105 0.439 ;
      RECT 4.091 0.738 4.105 0.793 ;
      RECT 4.000 0.738 4.091 0.819 ;
      RECT 4.059 0.323 4.085 0.404 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.696 0.167 3.787 0.257 ;
      RECT 3.601 0.202 3.696 0.257 ;
      RECT 3.659 0.683 3.680 0.764 ;
      RECT 3.601 0.567 3.659 0.764 ;
      RECT 3.589 0.202 3.601 0.764 ;
      RECT 3.557 0.202 3.589 0.633 ;
      RECT 3.540 0.202 3.557 0.621 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.057 0.335 1.191 0.494 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.213 0.512 0.329 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.352 -0.080 4.400 0.080 ;
      RECT 4.261 -0.080 4.352 0.122 ;
      RECT 4.000 -0.080 4.261 0.080 ;
      RECT 3.909 -0.080 4.000 0.122 ;
      RECT 3.573 -0.080 3.909 0.080 ;
      RECT 3.483 -0.080 3.573 0.122 ;
      RECT 3.051 -0.080 3.483 0.080 ;
      RECT 2.960 -0.080 3.051 0.287 ;
      RECT 2.353 -0.080 2.960 0.080 ;
      RECT 2.263 -0.080 2.353 0.329 ;
      RECT 1.776 -0.080 2.263 0.080 ;
      RECT 1.685 -0.080 1.776 0.287 ;
      RECT 0.837 -0.080 1.685 0.080 ;
      RECT 0.747 -0.080 0.837 0.122 ;
      RECT 0.323 -0.080 0.747 0.080 ;
      RECT 0.323 0.358 0.331 0.409 ;
      RECT 0.232 -0.080 0.323 0.409 ;
      RECT 0.000 -0.080 0.232 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.293 1.120 4.400 1.280 ;
      RECT 4.203 1.078 4.293 1.280 ;
      RECT 3.883 1.120 4.203 1.280 ;
      RECT 3.792 1.078 3.883 1.280 ;
      RECT 3.355 1.120 3.792 1.280 ;
      RECT 2.888 1.078 3.355 1.280 ;
      RECT 2.275 1.120 2.888 1.280 ;
      RECT 1.933 1.078 2.275 1.280 ;
      RECT 1.093 1.120 1.933 1.280 ;
      RECT 1.003 1.065 1.093 1.280 ;
      RECT 0.351 1.120 1.003 1.280 ;
      RECT 0.260 1.078 0.351 1.280 ;
      RECT 0.000 1.120 0.260 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.944 0.933 4.035 1.038 ;
      RECT 3.937 0.933 3.944 0.988 ;
      RECT 3.876 0.379 3.937 0.988 ;
      RECT 3.787 0.379 3.876 0.433 ;
      RECT 3.680 0.933 3.876 0.988 ;
      RECT 3.753 0.544 3.815 0.874 ;
      RECT 3.696 0.352 3.787 0.433 ;
      RECT 3.525 0.819 3.753 0.874 ;
      RECT 3.589 0.933 3.680 1.040 ;
      RECT 3.365 0.933 3.589 0.988 ;
      RECT 3.464 0.730 3.525 0.874 ;
      RECT 3.364 0.730 3.464 0.785 ;
      RECT 3.275 0.907 3.365 0.988 ;
      RECT 3.303 0.423 3.364 0.785 ;
      RECT 3.264 0.423 3.303 0.477 ;
      RECT 3.112 0.730 3.303 0.785 ;
      RECT 3.203 0.275 3.264 0.477 ;
      RECT 3.133 0.560 3.224 0.640 ;
      RECT 3.173 0.275 3.203 0.427 ;
      RECT 2.872 0.373 3.173 0.427 ;
      RECT 2.651 0.573 3.133 0.627 ;
      RECT 3.083 0.730 3.112 0.881 ;
      RECT 3.036 0.730 3.083 0.943 ;
      RECT 3.021 0.800 3.036 0.943 ;
      RECT 2.627 0.888 3.021 0.943 ;
      RECT 2.811 0.276 2.872 0.427 ;
      RECT 2.709 0.276 2.811 0.331 ;
      RECT 2.619 0.250 2.709 0.331 ;
      RECT 2.621 0.573 2.651 0.752 ;
      RECT 2.536 0.819 2.627 1.012 ;
      RECT 2.560 0.412 2.621 0.752 ;
      RECT 2.269 0.412 2.560 0.467 ;
      RECT 2.392 0.698 2.560 0.752 ;
      RECT 2.376 0.535 2.467 0.615 ;
      RECT 2.331 0.698 2.392 1.008 ;
      RECT 2.267 0.561 2.376 0.615 ;
      RECT 1.679 0.954 2.331 1.008 ;
      RECT 2.179 0.412 2.269 0.493 ;
      RECT 2.205 0.561 2.267 0.899 ;
      RECT 1.956 0.844 2.205 0.899 ;
      RECT 2.116 0.263 2.156 0.344 ;
      RECT 2.116 0.625 2.125 0.706 ;
      RECT 2.055 0.150 2.116 0.706 ;
      RECT 2.020 0.150 2.055 0.205 ;
      RECT 2.035 0.625 2.055 0.706 ;
      RECT 1.953 0.540 1.956 0.899 ;
      RECT 1.895 0.226 1.953 0.899 ;
      RECT 1.892 0.226 1.895 0.598 ;
      RECT 1.660 0.517 1.892 0.598 ;
      RECT 1.599 0.370 1.819 0.425 ;
      RECT 1.677 0.926 1.679 1.008 ;
      RECT 1.587 0.926 1.677 1.019 ;
      RECT 1.537 0.368 1.599 0.857 ;
      RECT 1.476 0.926 1.587 0.988 ;
      RECT 1.496 0.368 1.537 0.425 ;
      RECT 1.435 0.219 1.496 0.425 ;
      RECT 1.415 0.658 1.476 0.988 ;
      RECT 1.413 0.219 1.435 0.274 ;
      RECT 1.352 0.658 1.415 0.713 ;
      RECT 0.941 0.933 1.415 0.988 ;
      RECT 1.323 0.193 1.413 0.274 ;
      RECT 1.263 0.776 1.353 0.857 ;
      RECT 1.291 0.329 1.352 0.713 ;
      RECT 1.261 0.329 1.291 0.410 ;
      RECT 0.819 0.802 1.263 0.857 ;
      RECT 1.109 0.179 1.200 0.260 ;
      RECT 0.681 0.193 1.109 0.248 ;
      RECT 0.856 0.302 0.947 0.375 ;
      RECT 0.880 0.933 0.941 1.050 ;
      RECT 0.528 0.995 0.880 1.050 ;
      RECT 0.565 0.302 0.856 0.357 ;
      RECT 0.757 0.802 0.819 0.936 ;
      RECT 0.612 0.881 0.757 0.936 ;
      RECT 0.605 0.724 0.696 0.805 ;
      RECT 0.620 0.154 0.681 0.248 ;
      RECT 0.384 0.154 0.620 0.208 ;
      RECT 0.555 0.724 0.605 0.779 ;
      RECT 0.489 0.302 0.565 0.424 ;
      RECT 0.485 0.700 0.555 0.779 ;
      RECT 0.467 0.858 0.528 1.050 ;
      RECT 0.485 0.343 0.489 0.424 ;
      RECT 0.475 0.343 0.485 0.779 ;
      RECT 0.424 0.369 0.475 0.779 ;
      RECT 0.152 0.858 0.467 0.913 ;
      RECT 0.091 0.319 0.152 0.913 ;
      RECT 0.048 0.319 0.091 0.400 ;
      RECT 0.048 0.720 0.091 0.801 ;
  END
END SDFFX2

MACRO OR4X2
  CLASS CORE ;
  FOREIGN OR4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.997 0.182 1.061 1.010 ;
      RECT 0.942 0.182 0.997 0.375 ;
      RECT 0.953 0.700 0.997 1.010 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.728 0.700 0.878 0.767 ;
      RECT 0.664 0.552 0.728 0.767 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.406 0.527 0.556 0.633 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.167 0.364 0.264 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.433 0.151 0.567 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.646 -0.080 1.100 0.080 ;
      RECT 0.551 -0.080 0.646 0.122 ;
      RECT 0.144 -0.080 0.551 0.080 ;
      RECT 0.050 -0.080 0.144 0.122 ;
      RECT 0.000 -0.080 0.050 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.836 1.120 1.100 1.280 ;
      RECT 0.742 1.078 0.836 1.280 ;
      RECT 0.000 1.120 0.742 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.876 0.462 0.918 0.576 ;
      RECT 0.812 0.333 0.876 0.576 ;
      RECT 0.669 0.333 0.812 0.388 ;
      RECT 0.575 0.320 0.669 0.401 ;
      RECT 0.285 0.333 0.575 0.388 ;
      RECT 0.279 0.320 0.285 0.388 ;
      RECT 0.215 0.320 0.279 0.717 ;
      RECT 0.144 0.662 0.215 0.717 ;
      RECT 0.081 0.662 0.144 0.924 ;
      RECT 0.050 0.731 0.081 0.924 ;
  END
END OR4X2

MACRO OR3X2
  CLASS CORE ;
  FOREIGN OR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.039 0.182 1.061 0.500 ;
      RECT 0.975 0.182 1.039 1.010 ;
      RECT 0.956 0.182 0.975 0.500 ;
      RECT 0.944 0.705 0.975 1.010 ;
      RECT 0.944 0.182 0.956 0.375 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.586 0.601 0.700 0.775 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.506 0.423 0.539 0.507 ;
      RECT 0.411 0.423 0.506 0.518 ;
      RECT 0.383 0.423 0.411 0.507 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.186 0.567 0.322 0.668 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.839 -0.080 1.100 0.080 ;
      RECT 0.744 -0.080 0.839 0.211 ;
      RECT 0.375 -0.080 0.744 0.080 ;
      RECT 0.281 -0.080 0.375 0.122 ;
      RECT 0.000 -0.080 0.281 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.817 1.120 1.100 1.280 ;
      RECT 0.722 1.078 0.817 1.280 ;
      RECT 0.000 1.120 0.722 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.851 0.481 0.862 0.568 ;
      RECT 0.787 0.313 0.851 0.568 ;
      RECT 0.147 0.313 0.787 0.368 ;
      RECT 0.161 0.756 0.256 0.949 ;
      RECT 0.110 0.756 0.161 0.811 ;
      RECT 0.110 0.300 0.147 0.381 ;
      RECT 0.046 0.300 0.110 0.811 ;
  END
END OR3X2

MACRO OR2X2
  CLASS CORE ;
  FOREIGN OR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.589 0.196 0.650 0.914 ;
      RECT 0.548 0.196 0.589 0.389 ;
      RECT 0.546 0.721 0.589 0.914 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.414 0.337 0.558 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.393 0.138 0.544 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 -0.080 0.700 0.080 ;
      RECT 0.345 -0.080 0.435 0.122 ;
      RECT 0.138 -0.080 0.345 0.080 ;
      RECT 0.048 -0.080 0.138 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.435 1.120 0.700 1.280 ;
      RECT 0.345 1.078 0.435 1.280 ;
      RECT 0.000 1.120 0.345 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.460 0.502 0.528 0.583 ;
      RECT 0.399 0.279 0.460 0.776 ;
      RECT 0.286 0.279 0.399 0.333 ;
      RECT 0.138 0.721 0.399 0.776 ;
      RECT 0.196 0.252 0.286 0.333 ;
      RECT 0.048 0.721 0.138 0.802 ;
  END
END OR2X2

MACRO OAI33X2
  CLASS CORE ;
  FOREIGN OAI33X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.116 0.324 2.178 0.894 ;
      RECT 1.264 0.324 2.116 0.379 ;
      RECT 2.065 0.833 2.116 0.894 ;
      RECT 1.641 0.839 2.065 0.894 ;
      RECT 1.549 0.839 1.641 1.050 ;
      RECT 0.633 0.839 1.549 0.894 ;
      RECT 0.541 0.826 0.633 0.907 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.027 0.535 1.056 0.615 ;
      RECT 0.965 0.535 1.027 0.748 ;
      RECT 0.139 0.693 0.965 0.748 ;
      RECT 0.139 0.536 0.142 0.617 ;
      RECT 0.078 0.536 0.139 0.748 ;
      RECT 0.058 0.536 0.078 0.627 ;
      RECT 0.051 0.536 0.058 0.617 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.862 0.433 0.877 0.556 ;
      RECT 0.765 0.433 0.862 0.627 ;
      RECT 0.383 0.433 0.765 0.488 ;
      RECT 0.294 0.433 0.383 0.556 ;
      RECT 0.292 0.475 0.294 0.556 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.477 0.549 0.670 0.633 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.993 0.567 2.055 0.761 ;
      RECT 1.181 0.706 1.993 0.761 ;
      RECT 1.181 0.300 1.182 0.455 ;
      RECT 1.119 0.300 1.181 0.761 ;
      RECT 1.091 0.300 1.119 0.455 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.779 0.457 1.840 0.555 ;
      RECT 1.358 0.457 1.779 0.512 ;
      RECT 1.347 0.439 1.358 0.512 ;
      RECT 1.285 0.439 1.347 0.555 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.473 0.567 1.659 0.651 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.635 -0.080 2.300 0.080 ;
      RECT 0.544 -0.080 0.635 0.211 ;
      RECT 0.139 -0.080 0.544 0.080 ;
      RECT 0.048 -0.080 0.139 0.211 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.145 1.120 2.300 1.280 ;
      RECT 2.053 1.078 2.145 1.280 ;
      RECT 1.137 1.120 2.053 1.280 ;
      RECT 1.045 1.078 1.137 1.280 ;
      RECT 0.139 1.120 1.045 1.280 ;
      RECT 0.048 0.817 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.903 0.158 2.090 0.213 ;
      RECT 0.842 0.158 0.903 0.379 ;
      RECT 0.260 0.324 0.842 0.379 ;
  END
END OAI33X2

MACRO OAI32X2
  CLASS CORE ;
  FOREIGN OAI32X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.759 0.356 1.822 0.964 ;
      RECT 1.696 0.356 1.759 0.411 ;
      RECT 1.675 0.839 1.759 0.964 ;
      RECT 1.625 0.343 1.696 0.411 ;
      RECT 1.533 0.910 1.675 0.964 ;
      RECT 1.532 0.343 1.625 0.424 ;
      RECT 1.439 0.896 1.533 0.977 ;
      RECT 1.171 0.356 1.532 0.411 ;
      RECT 0.983 0.910 1.439 0.964 ;
      RECT 1.077 0.343 1.171 0.424 ;
      RECT 0.920 0.910 0.983 1.037 ;
      RECT 0.850 0.967 0.920 1.037 ;
      RECT 0.650 0.982 0.850 1.037 ;
      RECT 0.556 0.969 0.650 1.050 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.558 0.479 1.652 0.560 ;
      RECT 1.245 0.479 1.558 0.533 ;
      RECT 1.213 0.479 1.245 0.623 ;
      RECT 1.150 0.479 1.213 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.322 0.598 1.467 0.761 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.025 0.614 1.055 0.706 ;
      RECT 0.961 0.614 1.025 0.771 ;
      RECT 0.775 0.717 0.961 0.771 ;
      RECT 0.712 0.717 0.775 0.887 ;
      RECT 0.337 0.832 0.712 0.887 ;
      RECT 0.274 0.639 0.337 0.887 ;
      RECT 0.209 0.639 0.274 0.706 ;
      RECT 0.194 0.613 0.209 0.706 ;
      RECT 0.116 0.573 0.194 0.706 ;
      RECT 0.059 0.573 0.116 0.627 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.777 0.479 0.871 0.631 ;
      RECT 0.766 0.492 0.777 0.631 ;
      RECT 0.395 0.492 0.766 0.546 ;
      RECT 0.302 0.479 0.395 0.560 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.463 0.614 0.584 0.761 ;
      RECT 0.423 0.706 0.463 0.761 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.697 -0.080 2.000 0.080 ;
      RECT 0.603 -0.080 0.697 0.211 ;
      RECT 0.187 -0.080 0.603 0.080 ;
      RECT 0.094 -0.080 0.187 0.211 ;
      RECT 0.000 -0.080 0.094 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.897 1.120 2.000 1.280 ;
      RECT 1.803 1.078 1.897 1.280 ;
      RECT 1.169 1.120 1.803 1.280 ;
      RECT 1.076 1.078 1.169 1.280 ;
      RECT 0.143 1.120 1.076 1.280 ;
      RECT 0.050 0.877 0.143 1.280 ;
      RECT 0.000 1.120 0.050 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.227 0.150 1.450 0.231 ;
      RECT 0.931 0.163 1.227 0.218 ;
      RECT 0.868 0.163 0.931 0.424 ;
      RECT 0.837 0.343 0.868 0.424 ;
      RECT 0.493 0.356 0.837 0.411 ;
      RECT 0.270 0.343 0.493 0.424 ;
  END
END OAI32X2

MACRO OAI31X2
  CLASS CORE ;
  FOREIGN OAI31X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.339 0.343 1.368 0.439 ;
      RECT 1.216 0.804 1.343 0.911 ;
      RECT 1.277 0.343 1.339 0.512 ;
      RECT 1.216 0.457 1.277 0.512 ;
      RECT 1.154 0.457 1.216 0.911 ;
      RECT 1.125 0.839 1.154 0.911 ;
      RECT 0.636 0.856 1.125 0.911 ;
      RECT 0.544 0.856 0.636 1.049 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.282 0.567 1.399 0.719 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.037 0.614 1.083 0.695 ;
      RECT 0.991 0.614 1.037 0.792 ;
      RECT 0.975 0.627 0.991 0.792 ;
      RECT 0.947 0.706 0.975 0.792 ;
      RECT 0.236 0.737 0.947 0.792 ;
      RECT 0.205 0.700 0.236 0.792 ;
      RECT 0.143 0.614 0.205 0.792 ;
      RECT 0.113 0.614 0.143 0.695 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.873 0.539 0.902 0.620 ;
      RECT 0.811 0.445 0.873 0.620 ;
      RECT 0.475 0.445 0.811 0.500 ;
      RECT 0.413 0.439 0.475 0.500 ;
      RECT 0.393 0.445 0.413 0.500 ;
      RECT 0.331 0.445 0.393 0.620 ;
      RECT 0.294 0.539 0.331 0.620 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.479 0.567 0.673 0.668 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.024 -0.080 1.600 0.080 ;
      RECT 0.932 -0.080 1.024 0.122 ;
      RECT 0.646 -0.080 0.932 0.080 ;
      RECT 0.555 -0.080 0.646 0.122 ;
      RECT 0.291 -0.080 0.555 0.080 ;
      RECT 0.199 -0.080 0.291 0.122 ;
      RECT 0.000 -0.080 0.199 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.537 1.120 1.600 1.280 ;
      RECT 1.445 0.821 1.537 1.280 ;
      RECT 1.158 1.120 1.445 1.280 ;
      RECT 1.067 1.078 1.158 1.280 ;
      RECT 0.140 1.120 1.067 1.280 ;
      RECT 0.048 0.877 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.859 0.336 1.174 0.390 ;
      RECT 0.797 0.151 0.859 0.390 ;
      RECT 0.711 0.151 0.797 0.365 ;
      RECT 0.496 0.311 0.711 0.365 ;
      RECT 0.404 0.298 0.496 0.379 ;
      RECT 0.140 0.324 0.404 0.379 ;
      RECT 0.048 0.298 0.140 0.379 ;
  END
END OAI31X2

MACRO OAI2BB1X2
  CLASS CORE ;
  FOREIGN OAI2BB1X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.033 0.292 1.054 0.627 ;
      RECT 0.989 0.292 1.033 0.731 ;
      RECT 0.889 0.292 0.989 0.346 ;
      RECT 0.968 0.573 0.989 0.731 ;
      RECT 0.917 0.676 0.968 0.731 ;
      RECT 0.822 0.676 0.917 0.757 ;
      RECT 0.794 0.265 0.889 0.346 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.535 0.379 0.703 0.507 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.060 0.400 0.165 0.533 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.423 0.567 0.568 0.633 ;
      RECT 0.359 0.542 0.423 0.633 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.249 -0.080 1.300 0.080 ;
      RECT 1.154 -0.080 1.249 0.289 ;
      RECT 0.518 -0.080 1.154 0.080 ;
      RECT 0.422 -0.080 0.518 0.289 ;
      RECT 0.000 -0.080 0.422 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.109 1.120 1.300 1.280 ;
      RECT 1.013 1.078 1.109 1.280 ;
      RECT 0.737 1.120 1.013 1.280 ;
      RECT 0.642 0.972 0.737 1.280 ;
      RECT 0.298 1.120 0.642 1.280 ;
      RECT 0.203 1.078 0.298 1.280 ;
      RECT 0.000 1.120 0.203 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.833 0.468 0.864 0.549 ;
      RECT 0.768 0.468 0.833 0.621 ;
      RECT 0.756 0.567 0.768 0.621 ;
      RECT 0.691 0.567 0.756 0.823 ;
      RECT 0.523 0.768 0.691 0.823 ;
      RECT 0.428 0.768 0.523 0.849 ;
      RECT 0.294 0.768 0.428 0.823 ;
      RECT 0.229 0.280 0.294 0.823 ;
      RECT 0.146 0.280 0.229 0.335 ;
      RECT 0.051 0.254 0.146 0.335 ;
  END
END OAI2BB1X2

MACRO OAI22X2
  CLASS CORE ;
  FOREIGN OAI22X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.496 0.288 1.558 0.833 ;
      RECT 1.401 0.288 1.496 0.343 ;
      RECT 1.441 0.720 1.496 0.833 ;
      RECT 1.364 0.746 1.441 0.833 ;
      RECT 1.309 0.262 1.401 0.343 ;
      RECT 1.282 0.746 1.364 0.894 ;
      RECT 1.045 0.288 1.309 0.343 ;
      RECT 0.843 0.746 1.282 0.801 ;
      RECT 0.954 0.262 1.045 0.343 ;
      RECT 0.752 0.720 0.843 0.801 ;
      RECT 0.140 0.746 0.752 0.801 ;
      RECT 0.048 0.720 0.140 0.801 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.339 0.508 0.558 0.589 ;
      RECT 0.298 0.535 0.339 0.589 ;
      RECT 0.236 0.535 0.298 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.723 0.473 0.754 0.554 ;
      RECT 0.663 0.398 0.723 0.554 ;
      RECT 0.661 0.398 0.663 0.540 ;
      RECT 0.140 0.398 0.661 0.452 ;
      RECT 0.048 0.398 0.140 0.554 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.104 0.412 1.239 0.554 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.343 0.583 1.434 0.664 ;
      RECT 1.009 0.610 1.343 0.664 ;
      RECT 0.948 0.573 1.009 0.664 ;
      RECT 0.843 0.560 0.948 0.664 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.646 -0.080 1.600 0.080 ;
      RECT 0.555 -0.080 0.646 0.122 ;
      RECT 0.162 -0.080 0.555 0.080 ;
      RECT 0.070 -0.080 0.162 0.122 ;
      RECT 0.000 -0.080 0.070 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.188 1.120 1.600 1.280 ;
      RECT 1.096 0.911 1.188 1.280 ;
      RECT 0.496 1.120 1.096 1.280 ;
      RECT 0.404 0.911 0.496 1.280 ;
      RECT 0.000 1.120 0.404 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.760 0.261 0.851 0.342 ;
      RECT 0.496 0.287 0.760 0.342 ;
      RECT 0.404 0.261 0.496 0.342 ;
      RECT 0.140 0.287 0.404 0.342 ;
      RECT 0.048 0.261 0.140 0.342 ;
  END
END OAI22X2

MACRO OAI222X2
  CLASS CORE ;
  FOREIGN OAI222X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.274 0.331 2.335 0.888 ;
      RECT 1.861 0.331 2.274 0.386 ;
      RECT 2.197 0.833 2.274 0.888 ;
      RECT 2.136 0.833 2.197 0.894 ;
      RECT 1.964 0.839 2.136 0.894 ;
      RECT 1.849 0.839 1.964 0.920 ;
      RECT 1.271 0.839 1.849 0.894 ;
      RECT 1.154 0.839 1.271 0.920 ;
      RECT 0.588 0.839 1.154 0.894 ;
      RECT 0.499 0.839 0.588 0.920 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.185 0.675 2.214 0.730 ;
      RECT 2.125 0.675 2.185 0.743 ;
      RECT 1.733 0.688 2.125 0.743 ;
      RECT 1.673 0.573 1.733 0.743 ;
      RECT 1.616 0.573 1.673 0.627 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.943 0.498 2.043 0.633 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.290 0.552 0.827 0.607 ;
      RECT 0.242 0.552 0.290 0.627 ;
      RECT 0.152 0.546 0.242 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.637 0.662 0.651 0.743 ;
      RECT 0.576 0.662 0.637 0.761 ;
      RECT 0.436 0.662 0.576 0.743 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.422 0.562 1.535 0.617 ;
      RECT 1.362 0.552 1.422 0.617 ;
      RECT 1.051 0.552 1.362 0.607 ;
      RECT 0.990 0.552 1.051 0.640 ;
      RECT 0.961 0.560 0.990 0.640 ;
      RECT 0.923 0.573 0.961 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.297 0.700 1.341 0.767 ;
      RECT 1.208 0.662 1.297 0.767 ;
      RECT 1.129 0.700 1.208 0.767 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 2.600 0.080 ;
      RECT 0.762 -0.080 0.851 0.211 ;
      RECT 0.473 -0.080 0.762 0.080 ;
      RECT 0.383 -0.080 0.473 0.211 ;
      RECT 0.137 -0.080 0.383 0.080 ;
      RECT 0.047 -0.080 0.137 0.211 ;
      RECT 0.000 -0.080 0.047 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.280 1.120 2.600 1.280 ;
      RECT 2.190 0.984 2.280 1.280 ;
      RECT 1.597 1.120 2.190 1.280 ;
      RECT 1.507 0.984 1.597 1.280 ;
      RECT 0.924 1.120 1.507 1.280 ;
      RECT 0.835 0.984 0.924 1.280 ;
      RECT 0.252 1.120 0.835 1.280 ;
      RECT 0.163 0.984 0.252 1.280 ;
      RECT 0.000 1.120 0.163 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.746 0.193 2.487 0.248 ;
      RECT 1.686 0.158 1.746 0.327 ;
      RECT 0.945 0.158 1.686 0.213 ;
      RECT 1.203 0.302 1.572 0.357 ;
      RECT 1.114 0.302 1.203 0.399 ;
      RECT 0.662 0.302 1.114 0.357 ;
      RECT 0.633 0.212 0.662 0.357 ;
      RECT 0.573 0.212 0.633 0.373 ;
      RECT 0.305 0.318 0.573 0.373 ;
      RECT 0.215 0.318 0.305 0.399 ;
  END
END OAI222X2

MACRO OAI221X2
  CLASS CORE ;
  FOREIGN OAI221X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.976 0.345 2.032 0.830 ;
      RECT 1.970 0.318 1.976 0.830 ;
      RECT 1.914 0.318 1.970 0.440 ;
      RECT 1.732 0.775 1.970 0.830 ;
      RECT 1.716 0.775 1.732 0.839 ;
      RECT 1.654 0.775 1.716 0.904 ;
      RECT 1.624 0.823 1.654 0.904 ;
      RECT 1.169 0.839 1.624 0.894 ;
      RECT 1.078 0.839 1.169 0.920 ;
      RECT 1.003 0.839 1.078 0.900 ;
      RECT 0.483 0.839 1.003 0.894 ;
      RECT 0.391 0.839 0.483 0.920 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.647 0.567 1.903 0.633 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.204 0.552 0.740 0.607 ;
      RECT 0.113 0.546 0.204 0.627 ;
      RECT 0.058 0.573 0.113 0.627 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.473 0.662 0.547 0.743 ;
      RECT 0.411 0.662 0.473 0.761 ;
      RECT 0.327 0.662 0.411 0.743 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.319 0.562 1.512 0.617 ;
      RECT 1.257 0.552 1.319 0.617 ;
      RECT 1.004 0.552 1.257 0.607 ;
      RECT 0.954 0.552 1.004 0.627 ;
      RECT 0.942 0.552 0.954 0.640 ;
      RECT 0.863 0.560 0.942 0.640 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.196 0.700 1.240 0.767 ;
      RECT 1.104 0.662 1.196 0.767 ;
      RECT 1.024 0.700 1.104 0.767 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.869 -0.080 2.300 0.080 ;
      RECT 0.777 -0.080 0.869 0.211 ;
      RECT 0.483 -0.080 0.777 0.080 ;
      RECT 0.391 -0.080 0.483 0.211 ;
      RECT 0.139 -0.080 0.391 0.080 ;
      RECT 0.048 -0.080 0.139 0.211 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.909 1.120 2.300 1.280 ;
      RECT 1.817 0.900 1.909 1.280 ;
      RECT 1.512 1.120 1.817 1.280 ;
      RECT 1.421 0.984 1.512 1.280 ;
      RECT 0.826 1.120 1.421 1.280 ;
      RECT 0.734 0.984 0.826 1.280 ;
      RECT 0.139 1.120 0.734 1.280 ;
      RECT 0.048 0.929 0.139 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.783 0.193 2.162 0.248 ;
      RECT 1.721 0.158 1.783 0.327 ;
      RECT 0.965 0.158 1.721 0.213 ;
      RECT 1.228 0.302 1.604 0.357 ;
      RECT 1.137 0.302 1.228 0.399 ;
      RECT 0.676 0.302 1.137 0.357 ;
      RECT 0.646 0.217 0.676 0.357 ;
      RECT 0.584 0.217 0.646 0.373 ;
      RECT 0.311 0.318 0.584 0.373 ;
      RECT 0.220 0.318 0.311 0.399 ;
  END
END OAI221X2

MACRO OAI21X2
  CLASS CORE ;
  FOREIGN OAI21X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.283 0.311 1.343 0.920 ;
      RECT 1.282 0.311 1.283 0.946 ;
      RECT 1.114 0.311 1.282 0.365 ;
      RECT 1.151 0.865 1.282 0.946 ;
      RECT 0.838 0.865 1.151 0.920 ;
      RECT 1.053 0.263 1.114 0.365 ;
      RECT 1.023 0.263 1.053 0.344 ;
      RECT 0.748 0.865 0.838 0.946 ;
      RECT 0.138 0.865 0.748 0.920 ;
      RECT 0.048 0.865 0.138 0.946 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 0.551 1.179 0.632 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.614 0.562 0.695 ;
      RECT 0.473 0.614 0.488 0.707 ;
      RECT 0.407 0.614 0.473 0.761 ;
      RECT 0.323 0.614 0.407 0.707 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.711 0.605 0.740 0.686 ;
      RECT 0.650 0.460 0.711 0.686 ;
      RECT 0.232 0.460 0.650 0.514 ;
      RECT 0.119 0.433 0.232 0.514 ;
      RECT 0.118 0.439 0.119 0.514 ;
      RECT 0.057 0.439 0.118 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.732 -0.080 1.400 0.080 ;
      RECT 0.642 -0.080 0.732 0.280 ;
      RECT 0.339 -0.080 0.642 0.080 ;
      RECT 0.249 -0.080 0.339 0.122 ;
      RECT 0.000 -0.080 0.249 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.039 1.120 1.400 1.280 ;
      RECT 0.949 1.078 1.039 1.280 ;
      RECT 0.488 1.120 0.949 1.280 ;
      RECT 0.398 1.078 0.488 1.280 ;
      RECT 0.000 1.120 0.398 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.275 0.175 1.305 0.256 ;
      RECT 1.214 0.154 1.275 0.256 ;
      RECT 0.923 0.154 1.214 0.208 ;
      RECT 0.894 0.154 0.923 0.283 ;
      RECT 0.862 0.154 0.894 0.405 ;
      RECT 0.833 0.202 0.862 0.405 ;
      RECT 0.541 0.350 0.833 0.405 ;
      RECT 0.526 0.223 0.541 0.405 ;
      RECT 0.480 0.221 0.526 0.405 ;
      RECT 0.451 0.221 0.480 0.304 ;
      RECT 0.138 0.221 0.451 0.276 ;
      RECT 0.048 0.195 0.138 0.276 ;
  END
END OAI21X2

MACRO OAI211X2
  CLASS CORE ;
  FOREIGN OAI211X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.631 0.310 1.694 0.755 ;
      RECT 1.319 0.310 1.631 0.364 ;
      RECT 1.561 0.700 1.631 0.755 ;
      RECT 1.541 0.700 1.561 0.761 ;
      RECT 1.499 0.700 1.541 0.920 ;
      RECT 1.478 0.706 1.499 0.920 ;
      RECT 1.320 0.865 1.478 0.920 ;
      RECT 1.184 0.865 1.320 0.946 ;
      RECT 1.298 0.306 1.319 0.364 ;
      RECT 1.205 0.283 1.298 0.364 ;
      RECT 0.862 0.865 1.184 0.920 ;
      RECT 0.769 0.865 0.862 0.952 ;
      RECT 0.142 0.865 0.769 0.920 ;
      RECT 0.049 0.865 0.142 0.946 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.538 0.419 1.568 0.500 ;
      RECT 1.475 0.419 1.538 0.627 ;
      RECT 1.013 0.573 1.475 0.627 ;
      RECT 0.950 0.460 1.013 0.627 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.364 0.439 1.381 0.494 ;
      RECT 1.140 0.426 1.364 0.507 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.502 0.614 0.578 0.695 ;
      RECT 0.487 0.614 0.502 0.707 ;
      RECT 0.419 0.614 0.487 0.761 ;
      RECT 0.333 0.614 0.419 0.707 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.731 0.605 0.761 0.686 ;
      RECT 0.668 0.460 0.731 0.686 ;
      RECT 0.239 0.460 0.668 0.514 ;
      RECT 0.215 0.433 0.239 0.514 ;
      RECT 0.123 0.426 0.215 0.514 ;
      RECT 0.121 0.439 0.123 0.514 ;
      RECT 0.059 0.439 0.121 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.753 -0.080 1.800 0.080 ;
      RECT 0.660 -0.080 0.753 0.280 ;
      RECT 0.349 -0.080 0.660 0.080 ;
      RECT 0.256 -0.080 0.349 0.122 ;
      RECT 0.000 -0.080 0.256 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.069 1.120 1.800 1.280 ;
      RECT 0.976 1.078 1.069 1.280 ;
      RECT 0.502 1.120 0.976 1.280 ;
      RECT 0.409 1.078 0.502 1.280 ;
      RECT 0.000 1.120 0.409 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.555 0.171 1.647 0.252 ;
      RECT 0.949 0.174 1.555 0.229 ;
      RECT 0.919 0.174 0.949 0.283 ;
      RECT 0.886 0.174 0.919 0.405 ;
      RECT 0.856 0.202 0.886 0.405 ;
      RECT 0.556 0.350 0.856 0.405 ;
      RECT 0.541 0.223 0.556 0.405 ;
      RECT 0.494 0.221 0.541 0.405 ;
      RECT 0.464 0.221 0.494 0.304 ;
      RECT 0.142 0.221 0.464 0.276 ;
      RECT 0.049 0.195 0.142 0.276 ;
  END
END OAI211X2

MACRO NOR4BBX2
  CLASS CORE ;
  FOREIGN NOR4BBX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.901 0.150 1.964 0.986 ;
      RECT 1.295 0.150 1.901 0.205 ;
      RECT 1.857 0.894 1.901 0.986 ;
      RECT 1.032 0.931 1.857 0.986 ;
      RECT 1.231 0.150 1.295 0.246 ;
      RECT 0.959 0.192 1.231 0.246 ;
      RECT 0.968 0.931 1.032 1.027 ;
      RECT 0.917 0.931 0.968 1.012 ;
      RECT 0.865 0.165 0.959 0.246 ;
      RECT 0.540 0.192 0.865 0.246 ;
      RECT 0.446 0.165 0.540 0.246 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.563 0.570 1.602 0.625 ;
      RECT 1.500 0.570 1.563 0.876 ;
      RECT 0.486 0.821 1.500 0.876 ;
      RECT 0.423 0.821 0.486 0.894 ;
      RECT 0.379 0.821 0.423 0.876 ;
      RECT 0.315 0.557 0.379 0.876 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.379 0.570 1.416 0.625 ;
      RECT 1.379 0.704 1.395 0.761 ;
      RECT 1.332 0.570 1.379 0.761 ;
      RECT 1.315 0.570 1.332 0.758 ;
      RECT 0.595 0.704 1.315 0.758 ;
      RECT 0.517 0.457 0.595 0.758 ;
      RECT 0.501 0.457 0.517 0.538 ;
     END
  END C

  PIN BN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.556 0.277 1.780 0.396 ;
     END
  END BN

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.249 0.433 0.348 0.500 ;
      RECT 0.160 0.380 0.249 0.500 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.168 -0.080 2.000 0.080 ;
      RECT 1.074 -0.080 1.168 0.122 ;
      RECT 0.749 -0.080 1.074 0.080 ;
      RECT 0.656 -0.080 0.749 0.122 ;
      RECT 0.342 -0.080 0.656 0.080 ;
      RECT 0.248 -0.080 0.342 0.198 ;
      RECT 0.000 -0.080 0.248 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.683 1.120 2.000 1.280 ;
      RECT 1.590 1.078 1.683 1.280 ;
      RECT 0.298 1.120 1.590 1.280 ;
      RECT 0.204 1.078 0.298 1.280 ;
      RECT 0.000 1.120 0.204 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.774 0.457 1.837 0.764 ;
      RECT 1.421 0.457 1.774 0.512 ;
      RECT 1.421 0.262 1.493 0.317 ;
      RECT 1.358 0.262 1.421 0.512 ;
      RECT 1.231 0.457 1.358 0.512 ;
      RECT 1.201 0.457 1.231 0.538 ;
      RECT 1.138 0.457 1.201 0.649 ;
      RECT 0.791 0.594 1.138 0.649 ;
      RECT 0.982 0.457 1.012 0.538 ;
      RECT 0.919 0.324 0.982 0.538 ;
      RECT 0.382 0.324 0.919 0.379 ;
      RECT 0.727 0.457 0.791 0.649 ;
      RECT 0.697 0.457 0.727 0.538 ;
      RECT 0.318 0.269 0.382 0.379 ;
      RECT 0.143 0.269 0.318 0.324 ;
      RECT 0.096 0.217 0.143 0.324 ;
      RECT 0.096 0.683 0.143 0.876 ;
      RECT 0.033 0.217 0.096 0.876 ;
  END
END NOR4BBX2

MACRO NOR4BX2
  CLASS CORE ;
  FOREIGN NOR4BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.675 0.192 1.737 0.894 ;
      RECT 1.658 0.192 1.675 0.306 ;
      RECT 1.140 0.839 1.675 0.894 ;
      RECT 0.949 0.192 1.658 0.246 ;
      RECT 1.058 0.833 1.140 0.900 ;
      RECT 0.965 0.826 1.058 0.907 ;
      RECT 0.856 0.179 0.949 0.260 ;
      RECT 0.442 0.192 0.856 0.246 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.580 0.557 1.612 0.638 ;
      RECT 1.519 0.557 1.580 0.761 ;
      RECT 1.518 0.570 1.519 0.761 ;
      RECT 0.419 0.706 1.518 0.761 ;
      RECT 0.390 0.700 0.419 0.761 ;
      RECT 0.297 0.569 0.390 0.761 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.396 1.561 0.500 ;
      RECT 1.400 0.343 1.480 0.500 ;
      RECT 0.682 0.343 1.400 0.398 ;
      RECT 0.641 0.343 0.682 0.439 ;
      RECT 0.578 0.343 0.641 0.533 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.139 0.452 1.276 0.627 ;
      RECT 0.840 0.452 1.139 0.507 ;
      RECT 0.747 0.452 0.840 0.533 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.222 0.433 0.322 0.513 ;
      RECT 0.160 0.395 0.222 0.513 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.156 -0.080 1.800 0.080 ;
      RECT 1.064 -0.080 1.156 0.122 ;
      RECT 0.742 -0.080 1.064 0.080 ;
      RECT 0.649 -0.080 0.742 0.122 ;
      RECT 0.338 -0.080 0.649 0.080 ;
      RECT 0.245 -0.080 0.338 0.198 ;
      RECT 0.000 -0.080 0.245 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.724 1.120 1.800 1.280 ;
      RECT 1.631 1.078 1.724 1.280 ;
      RECT 0.327 1.120 1.631 1.280 ;
      RECT 0.235 1.078 0.327 1.280 ;
      RECT 0.000 1.120 0.235 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.926 0.570 1.023 0.643 ;
      RECT 0.515 0.588 0.926 0.643 ;
      RECT 0.453 0.301 0.515 0.643 ;
      RECT 0.359 0.301 0.453 0.356 ;
      RECT 0.296 0.268 0.359 0.356 ;
      RECT 0.142 0.268 0.296 0.323 ;
      RECT 0.097 0.217 0.142 0.323 ;
      RECT 0.097 0.683 0.142 0.876 ;
      RECT 0.034 0.217 0.097 0.876 ;
  END
END NOR4BX2

MACRO NOR4X2
  CLASS CORE ;
  FOREIGN NOR4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.287 1.542 1.008 ;
      RECT 0.813 0.287 1.480 0.342 ;
      RECT 1.460 0.894 1.480 1.008 ;
      RECT 0.853 0.954 1.460 1.008 ;
      RECT 0.761 0.954 0.853 1.035 ;
      RECT 0.722 0.261 0.813 0.342 ;
      RECT 0.338 0.287 0.722 0.342 ;
      RECT 0.246 0.261 0.338 0.342 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.387 0.556 1.417 0.637 ;
      RECT 1.325 0.556 1.387 0.899 ;
      RECT 0.238 0.844 1.325 0.899 ;
      RECT 0.176 0.556 0.238 0.899 ;
      RECT 0.055 0.556 0.176 0.637 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.174 0.396 1.236 0.789 ;
      RECT 1.145 0.396 1.174 0.477 ;
      RECT 0.475 0.735 1.174 0.789 ;
      RECT 0.427 0.706 0.475 0.789 ;
      RECT 0.365 0.556 0.427 0.789 ;
      RECT 0.335 0.556 0.365 0.637 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.069 0.556 1.099 0.637 ;
      RECT 1.007 0.444 1.069 0.637 ;
      RECT 0.653 0.444 1.007 0.499 ;
      RECT 0.607 0.439 0.653 0.499 ;
      RECT 0.517 0.439 0.607 0.538 ;
      RECT 0.516 0.457 0.517 0.538 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.710 0.555 0.878 0.636 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.018 -0.080 1.600 0.080 ;
      RECT 0.927 -0.080 1.018 0.122 ;
      RECT 0.593 -0.080 0.927 0.080 ;
      RECT 0.501 -0.080 0.593 0.122 ;
      RECT 0.140 -0.080 0.501 0.080 ;
      RECT 0.048 -0.080 0.140 0.225 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.534 1.120 1.600 1.280 ;
      RECT 1.442 1.078 1.534 1.280 ;
      RECT 0.140 1.120 1.442 1.280 ;
      RECT 0.048 1.078 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
END NOR4X2

MACRO NOR3BX2
  CLASS CORE ;
  FOREIGN NOR3BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.270 0.192 1.331 0.861 ;
      RECT 1.262 0.192 1.270 0.306 ;
      RECT 1.262 0.761 1.270 0.861 ;
      RECT 0.973 0.192 1.262 0.246 ;
      RECT 0.993 0.806 1.262 0.861 ;
      RECT 0.932 0.806 0.993 0.894 ;
      RECT 0.883 0.165 0.973 0.246 ;
      RECT 0.843 0.806 0.932 0.861 ;
      RECT 0.570 0.192 0.883 0.246 ;
      RECT 0.753 0.806 0.843 0.895 ;
      RECT 0.480 0.165 0.570 0.246 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.180 0.394 1.209 0.475 ;
      RECT 1.119 0.324 1.180 0.475 ;
      RECT 0.467 0.324 1.119 0.379 ;
      RECT 0.467 0.573 0.468 0.627 ;
      RECT 0.406 0.324 0.467 0.627 ;
      RECT 0.387 0.494 0.406 0.627 ;
      RECT 0.365 0.536 0.387 0.627 ;
      RECT 0.335 0.536 0.365 0.617 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.057 0.555 1.086 0.636 ;
      RECT 0.996 0.461 1.057 0.636 ;
      RECT 0.643 0.461 0.996 0.515 ;
      RECT 0.619 0.439 0.643 0.515 ;
      RECT 0.558 0.439 0.619 0.542 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.273 0.306 0.293 0.361 ;
      RECT 0.212 0.306 0.273 0.457 ;
      RECT 0.174 0.376 0.212 0.457 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.772 -0.080 1.400 0.080 ;
      RECT 0.681 -0.080 0.772 0.122 ;
      RECT 0.379 -0.080 0.681 0.080 ;
      RECT 0.289 -0.080 0.379 0.198 ;
      RECT 0.000 -0.080 0.289 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 1.120 1.400 1.280 ;
      RECT 1.246 0.932 1.336 1.280 ;
      RECT 0.345 1.120 1.246 1.280 ;
      RECT 0.255 0.897 0.345 1.280 ;
      RECT 0.000 1.120 0.255 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.846 0.570 0.875 0.625 ;
      RECT 0.785 0.570 0.846 0.751 ;
      RECT 0.138 0.696 0.785 0.751 ;
      RECT 0.109 0.198 0.151 0.282 ;
      RECT 0.109 0.670 0.138 0.751 ;
      RECT 0.048 0.198 0.109 0.751 ;
  END
END NOR3BX2

MACRO NOR3X2
  CLASS CORE ;
  FOREIGN NOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.175 0.255 1.240 0.855 ;
      RECT 0.754 0.255 1.175 0.310 ;
      RECT 1.154 0.767 1.175 0.855 ;
      RECT 0.687 0.800 1.154 0.855 ;
      RECT 0.658 0.151 0.754 0.344 ;
      RECT 0.591 0.800 0.687 0.890 ;
      RECT 0.349 0.289 0.658 0.344 ;
      RECT 0.253 0.151 0.349 0.344 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.007 0.537 1.088 0.744 ;
      RECT 0.214 0.689 1.007 0.744 ;
      RECT 0.149 0.573 0.214 0.744 ;
      RECT 0.118 0.573 0.149 0.707 ;
      RECT 0.058 0.573 0.118 0.627 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.913 0.377 0.943 0.458 ;
      RECT 0.848 0.377 0.913 0.635 ;
      RECT 0.847 0.377 0.848 0.458 ;
      RECT 0.416 0.580 0.848 0.635 ;
      RECT 0.415 0.458 0.416 0.635 ;
      RECT 0.352 0.445 0.415 0.635 ;
      RECT 0.321 0.445 0.352 0.539 ;
      RECT 0.311 0.445 0.321 0.500 ;
      RECT 0.246 0.439 0.311 0.500 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.498 0.439 0.682 0.525 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.552 -0.080 1.300 0.080 ;
      RECT 0.456 -0.080 0.552 0.211 ;
      RECT 0.146 -0.080 0.456 0.080 ;
      RECT 0.051 -0.080 0.146 0.211 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.204 1.120 1.300 1.280 ;
      RECT 1.109 0.925 1.204 1.280 ;
      RECT 0.146 1.120 1.109 1.280 ;
      RECT 0.051 0.876 0.146 1.280 ;
      RECT 0.000 1.120 0.051 1.280 ;
     END
  END VDD
END NOR3X2

MACRO NOR2BX2
  CLASS CORE ;
  FOREIGN NOR2BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.997 0.308 1.061 0.767 ;
      RECT 0.850 0.308 0.997 0.363 ;
      RECT 0.976 0.706 0.997 0.767 ;
      RECT 0.689 0.712 0.976 0.767 ;
      RECT 0.756 0.282 0.850 0.363 ;
      RECT 0.594 0.712 0.689 0.793 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.847 0.418 0.928 0.565 ;
      RECT 0.511 0.418 0.847 0.473 ;
      RECT 0.436 0.300 0.511 0.473 ;
      RECT 0.406 0.300 0.436 0.514 ;
      RECT 0.357 0.418 0.406 0.514 ;
      RECT 0.342 0.433 0.357 0.514 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.050 0.457 0.144 0.633 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 -0.080 1.100 0.080 ;
      RECT 0.956 -0.080 1.050 0.228 ;
      RECT 0.636 -0.080 0.956 0.080 ;
      RECT 0.542 -0.080 0.636 0.122 ;
      RECT 0.000 -0.080 0.542 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 1.120 1.100 1.280 ;
      RECT 0.956 1.078 1.050 1.280 ;
      RECT 0.322 1.120 0.956 1.280 ;
      RECT 0.228 1.078 0.322 1.280 ;
      RECT 0.000 1.120 0.228 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.622 0.538 0.717 0.626 ;
      RECT 0.272 0.571 0.622 0.626 ;
      RECT 0.208 0.312 0.272 0.802 ;
      RECT 0.144 0.312 0.208 0.367 ;
      RECT 0.144 0.748 0.208 0.802 ;
      RECT 0.050 0.286 0.144 0.367 ;
      RECT 0.050 0.748 0.144 0.829 ;
  END
END NOR2BX2

MACRO NOR2X2
  CLASS CORE ;
  FOREIGN NOR2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.862 0.308 0.867 0.761 ;
      RECT 0.805 0.308 0.862 0.767 ;
      RECT 0.655 0.308 0.805 0.363 ;
      RECT 0.779 0.706 0.805 0.767 ;
      RECT 0.496 0.712 0.779 0.767 ;
      RECT 0.562 0.170 0.655 0.363 ;
      RECT 0.404 0.712 0.496 0.793 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.652 0.418 0.742 0.564 ;
      RECT 0.229 0.418 0.652 0.473 ;
      RECT 0.120 0.418 0.229 0.518 ;
      RECT 0.059 0.418 0.120 0.494 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.327 0.538 0.502 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.228 ;
      RECT 0.458 -0.080 0.758 0.080 ;
      RECT 0.365 -0.080 0.458 0.340 ;
      RECT 0.000 -0.080 0.365 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.758 1.078 0.851 1.280 ;
      RECT 0.142 1.120 0.758 1.280 ;
      RECT 0.049 1.078 0.142 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
END NOR2X2

MACRO NAND4BBX2
  CLASS CORE ;
  FOREIGN NAND4BBX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.884 0.195 1.961 0.973 ;
      RECT 0.990 0.195 1.884 0.262 ;
      RECT 1.879 0.573 1.884 0.973 ;
      RECT 1.868 0.573 1.879 0.644 ;
      RECT 1.857 0.893 1.879 0.973 ;
      RECT 1.055 0.901 1.857 0.973 ;
      RECT 0.972 0.870 1.055 0.973 ;
      RECT 0.897 0.150 0.990 0.343 ;
      RECT 0.444 0.870 0.972 0.942 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.371 0.761 1.464 0.842 ;
      RECT 0.486 0.761 1.371 0.815 ;
      RECT 0.428 0.706 0.486 0.815 ;
      RECT 0.365 0.519 0.428 0.815 ;
      RECT 0.340 0.519 0.365 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.380 0.573 1.395 0.627 ;
      RECT 1.350 0.519 1.380 0.627 ;
      RECT 1.287 0.519 1.350 0.706 ;
      RECT 0.634 0.651 1.287 0.706 ;
      RECT 0.570 0.519 0.634 0.706 ;
      RECT 0.522 0.519 0.570 0.600 ;
     END
  END C

  PIN BN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.657 0.498 1.780 0.633 ;
     END
  END BN

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.043 0.433 0.147 0.574 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.663 -0.080 2.000 0.080 ;
      RECT 1.569 -0.080 1.663 0.122 ;
      RECT 0.318 -0.080 1.569 0.080 ;
      RECT 0.092 -0.080 0.318 0.122 ;
      RECT 0.000 -0.080 0.092 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.882 1.120 2.000 1.280 ;
      RECT 1.737 1.078 1.882 1.280 ;
      RECT 1.140 1.120 1.737 1.280 ;
      RECT 1.017 1.078 1.140 1.280 ;
      RECT 0.733 1.120 1.017 1.280 ;
      RECT 0.639 1.078 0.733 1.280 ;
      RECT 0.342 1.120 0.639 1.280 ;
      RECT 0.248 1.078 0.342 1.280 ;
      RECT 0.000 1.120 0.248 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.758 0.317 1.821 0.398 ;
      RECT 1.591 0.330 1.758 0.398 ;
      RECT 1.591 0.761 1.621 0.842 ;
      RECT 1.528 0.330 1.591 0.842 ;
      RECT 1.200 0.401 1.528 0.456 ;
      RECT 1.136 0.401 1.200 0.596 ;
      RECT 1.096 0.514 1.136 0.596 ;
      RECT 0.809 0.542 1.096 0.596 ;
      RECT 0.895 0.400 0.999 0.487 ;
      RECT 0.274 0.400 0.895 0.455 ;
      RECT 0.705 0.515 0.809 0.596 ;
      RECT 0.211 0.302 0.274 0.730 ;
      RECT 0.143 0.302 0.211 0.357 ;
      RECT 0.143 0.675 0.211 0.730 ;
      RECT 0.050 0.276 0.143 0.357 ;
      RECT 0.050 0.675 0.143 0.868 ;
  END
END NAND4BBX2

MACRO NAND4BX2
  CLASS CORE ;
  FOREIGN NAND4BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.800 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.740 0.195 1.741 0.633 ;
      RECT 1.665 0.195 1.740 0.973 ;
      RECT 1.658 0.195 1.665 0.306 ;
      RECT 1.658 0.564 1.665 0.973 ;
      RECT 0.987 0.195 1.658 0.262 ;
      RECT 1.045 0.901 1.658 0.973 ;
      RECT 0.963 0.870 1.045 0.973 ;
      RECT 0.895 0.150 0.987 0.343 ;
      RECT 0.439 0.870 0.963 0.942 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.357 0.761 1.450 0.842 ;
      RECT 0.481 0.761 1.357 0.815 ;
      RECT 0.424 0.706 0.481 0.815 ;
      RECT 0.419 0.519 0.424 0.815 ;
      RECT 0.361 0.519 0.419 0.761 ;
      RECT 0.340 0.519 0.361 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.377 0.573 1.381 0.627 ;
      RECT 1.347 0.519 1.377 0.627 ;
      RECT 1.285 0.519 1.347 0.706 ;
      RECT 0.627 0.651 1.285 0.706 ;
      RECT 0.565 0.519 0.627 0.706 ;
      RECT 0.521 0.519 0.565 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.188 0.439 1.201 0.494 ;
      RECT 1.118 0.433 1.188 0.596 ;
      RECT 1.085 0.514 1.118 0.596 ;
      RECT 0.800 0.542 1.085 0.596 ;
      RECT 0.698 0.515 0.800 0.596 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.042 0.433 0.146 0.574 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.653 -0.080 1.800 0.080 ;
      RECT 1.560 -0.080 1.653 0.122 ;
      RECT 0.322 -0.080 1.560 0.080 ;
      RECT 0.229 -0.080 0.322 0.122 ;
      RECT 0.000 -0.080 0.229 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.129 1.120 1.800 1.280 ;
      RECT 1.006 1.078 1.129 1.280 ;
      RECT 0.725 1.120 1.006 1.280 ;
      RECT 0.633 1.078 0.725 1.280 ;
      RECT 0.338 1.120 0.633 1.280 ;
      RECT 0.323 1.078 0.338 1.280 ;
      RECT 0.260 1.065 0.323 1.280 ;
      RECT 0.245 1.078 0.260 1.280 ;
      RECT 0.000 1.120 0.245 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.886 0.400 0.989 0.487 ;
      RECT 0.274 0.400 0.886 0.455 ;
      RECT 0.211 0.302 0.274 0.799 ;
      RECT 0.142 0.302 0.211 0.357 ;
      RECT 0.142 0.744 0.211 0.799 ;
      RECT 0.049 0.276 0.142 0.357 ;
      RECT 0.049 0.731 0.142 0.812 ;
  END
END NAND4BX2

MACRO NAND4X2
  CLASS CORE ;
  FOREIGN NAND4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 0.195 1.542 0.633 ;
      RECT 1.467 0.195 1.541 0.973 ;
      RECT 1.460 0.195 1.467 0.306 ;
      RECT 1.460 0.564 1.467 0.973 ;
      RECT 0.797 0.195 1.460 0.262 ;
      RECT 0.854 0.901 1.460 0.973 ;
      RECT 0.773 0.870 0.854 0.973 ;
      RECT 0.706 0.150 0.797 0.343 ;
      RECT 0.256 0.870 0.773 0.942 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.162 0.761 1.254 0.842 ;
      RECT 0.298 0.761 1.162 0.815 ;
      RECT 0.241 0.706 0.298 0.815 ;
      RECT 0.236 0.519 0.241 0.815 ;
      RECT 0.179 0.519 0.236 0.761 ;
      RECT 0.149 0.519 0.179 0.600 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.187 0.519 1.193 0.600 ;
      RECT 1.164 0.519 1.187 0.627 ;
      RECT 1.102 0.519 1.164 0.706 ;
      RECT 0.442 0.651 1.102 0.706 ;
      RECT 0.380 0.519 0.442 0.706 ;
      RECT 0.333 0.519 0.380 0.600 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.916 0.439 1.017 0.596 ;
      RECT 0.613 0.542 0.916 0.596 ;
      RECT 0.512 0.515 0.613 0.596 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.698 0.401 0.799 0.487 ;
      RECT 0.496 0.401 0.698 0.456 ;
      RECT 0.434 0.306 0.496 0.456 ;
      RECT 0.413 0.306 0.434 0.361 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.455 -0.080 1.600 0.080 ;
      RECT 1.363 -0.080 1.455 0.122 ;
      RECT 0.140 -0.080 1.363 0.080 ;
      RECT 0.048 -0.080 0.140 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.937 1.120 1.600 1.280 ;
      RECT 0.816 1.078 0.937 1.280 ;
      RECT 0.539 1.120 0.816 1.280 ;
      RECT 0.447 1.078 0.539 1.280 ;
      RECT 0.156 1.120 0.447 1.280 ;
      RECT 0.065 1.078 0.156 1.280 ;
      RECT 0.000 1.120 0.065 1.280 ;
     END
  END VDD
END NAND4X2

MACRO NAND3BX2
  CLASS CORE ;
  FOREIGN NAND3BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.651 0.689 0.741 0.770 ;
      RECT 0.567 0.164 0.658 0.245 ;
      RECT 0.643 0.689 0.651 0.767 ;
      RECT 0.407 0.700 0.643 0.767 ;
      RECT 0.294 0.177 0.567 0.232 ;
      RECT 0.373 0.689 0.407 0.767 ;
      RECT 0.294 0.689 0.373 0.770 ;
      RECT 0.282 0.177 0.294 0.770 ;
      RECT 0.233 0.177 0.282 0.767 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.033 0.462 1.047 0.543 ;
      RECT 0.972 0.462 1.033 0.881 ;
      RECT 0.957 0.462 0.972 0.543 ;
      RECT 0.172 0.826 0.972 0.881 ;
      RECT 0.111 0.439 0.172 0.881 ;
      RECT 0.082 0.439 0.111 0.573 ;
      RECT 0.057 0.439 0.082 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.838 0.507 0.870 0.588 ;
      RECT 0.737 0.433 0.838 0.604 ;
      RECT 0.445 0.549 0.737 0.604 ;
      RECT 0.355 0.514 0.445 0.604 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.358 0.467 1.363 0.594 ;
      RECT 1.267 0.433 1.358 0.594 ;
      RECT 1.262 0.467 1.267 0.594 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.161 -0.080 1.400 0.080 ;
      RECT 1.145 -0.080 1.161 0.122 ;
      RECT 1.055 -0.080 1.145 0.247 ;
      RECT 0.154 -0.080 1.055 0.080 ;
      RECT 0.064 -0.080 0.154 0.247 ;
      RECT 0.000 -0.080 0.064 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.148 1.120 1.400 1.280 ;
      RECT 1.058 0.952 1.148 1.280 ;
      RECT 0.561 1.120 1.058 1.280 ;
      RECT 0.471 0.952 0.561 1.280 ;
      RECT 0.192 1.120 0.471 1.280 ;
      RECT 0.102 0.952 0.192 1.280 ;
      RECT 0.000 1.120 0.102 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.262 0.279 1.352 0.379 ;
      RECT 1.262 0.702 1.352 0.783 ;
      RECT 1.201 0.324 1.262 0.379 ;
      RECT 1.201 0.702 1.262 0.757 ;
      RECT 1.140 0.324 1.201 0.757 ;
      RECT 0.658 0.324 1.140 0.379 ;
      RECT 0.597 0.324 0.658 0.490 ;
      RECT 0.567 0.410 0.597 0.490 ;
  END
END NAND3BX2

MACRO NAND3X2
  CLASS CORE ;
  FOREIGN NAND3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.691 0.689 0.786 0.770 ;
      RECT 0.602 0.164 0.698 0.245 ;
      RECT 0.682 0.689 0.691 0.761 ;
      RECT 0.518 0.706 0.682 0.761 ;
      RECT 0.312 0.190 0.602 0.245 ;
      RECT 0.432 0.700 0.518 0.770 ;
      RECT 0.312 0.689 0.432 0.770 ;
      RECT 0.300 0.190 0.312 0.770 ;
      RECT 0.248 0.190 0.300 0.761 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.096 0.573 1.111 0.706 ;
      RECT 1.031 0.573 1.096 0.881 ;
      RECT 1.016 0.573 1.031 0.706 ;
      RECT 0.183 0.826 1.031 0.881 ;
      RECT 0.167 0.460 0.183 0.881 ;
      RECT 0.118 0.439 0.167 0.881 ;
      RECT 0.087 0.439 0.118 0.573 ;
      RECT 0.060 0.439 0.087 0.494 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.907 0.493 0.923 0.588 ;
      RECT 0.868 0.433 0.907 0.588 ;
      RECT 0.782 0.433 0.868 0.604 ;
      RECT 0.473 0.549 0.782 0.604 ;
      RECT 0.377 0.514 0.473 0.604 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.602 0.300 0.698 0.490 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.232 -0.080 1.300 0.080 ;
      RECT 1.137 -0.080 1.232 0.122 ;
      RECT 0.163 -0.080 1.137 0.080 ;
      RECT 0.068 -0.080 0.163 0.122 ;
      RECT 0.000 -0.080 0.068 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.595 1.120 1.300 1.280 ;
      RECT 0.499 0.952 0.595 1.280 ;
      RECT 0.204 1.120 0.499 1.280 ;
      RECT 0.108 0.952 0.204 1.280 ;
      RECT 0.000 1.120 0.108 1.280 ;
     END
  END VDD
END NAND3X2

MACRO NAND2BX2
  CLASS CORE ;
  FOREIGN NAND2BX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.003 0.402 1.067 0.870 ;
      RECT 0.894 0.800 1.003 0.870 ;
      RECT 0.800 0.790 0.894 0.871 ;
      RECT 0.772 0.800 0.800 0.870 ;
      RECT 0.610 0.815 0.772 0.870 ;
      RECT 0.539 0.802 0.610 0.870 ;
      RECT 0.444 0.802 0.539 0.883 ;
      RECT 0.878 0.402 1.003 0.457 ;
      RECT 0.876 0.361 0.878 0.457 ;
      RECT 0.812 0.317 0.876 0.457 ;
      RECT 0.694 0.317 0.812 0.371 ;
      RECT 0.600 0.290 0.694 0.371 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.853 0.599 0.939 0.686 ;
      RECT 0.467 0.623 0.853 0.677 ;
      RECT 0.372 0.610 0.467 0.690 ;
     END
  END B

  PIN AN
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.047 0.452 0.142 0.627 ;
     END
  END AN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 -0.080 1.100 0.080 ;
      RECT 0.956 -0.080 1.050 0.278 ;
      RECT 0.328 -0.080 0.956 0.080 ;
      RECT 0.233 -0.080 0.328 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.050 1.120 1.100 1.280 ;
      RECT 0.353 1.078 1.050 1.280 ;
      RECT 0.000 1.120 0.353 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.639 0.433 0.733 0.514 ;
      RECT 0.272 0.446 0.639 0.501 ;
      RECT 0.208 0.311 0.272 0.757 ;
      RECT 0.144 0.311 0.208 0.368 ;
      RECT 0.144 0.702 0.208 0.757 ;
      RECT 0.050 0.279 0.144 0.368 ;
      RECT 0.050 0.702 0.144 0.783 ;
      RECT 0.049 0.292 0.050 0.368 ;
  END
END NAND2BX2

MACRO NAND2X2
  CLASS CORE ;
  FOREIGN NAND2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.795 0.402 0.858 0.770 ;
      RECT 0.680 0.402 0.795 0.457 ;
      RECT 0.779 0.704 0.795 0.770 ;
      RECT 0.251 0.704 0.779 0.758 ;
      RECT 0.618 0.249 0.680 0.457 ;
      RECT 0.599 0.249 0.618 0.306 ;
      RECT 0.502 0.249 0.599 0.304 ;
      RECT 0.409 0.223 0.502 0.304 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.668 0.558 0.731 0.645 ;
      RECT 0.301 0.577 0.668 0.632 ;
      RECT 0.200 0.573 0.301 0.632 ;
      RECT 0.185 0.573 0.200 0.627 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.398 0.400 0.551 0.520 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 -0.080 0.900 0.080 ;
      RECT 0.758 -0.080 0.851 0.289 ;
      RECT 0.142 -0.080 0.758 0.080 ;
      RECT 0.049 -0.080 0.142 0.122 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 1.120 0.900 1.280 ;
      RECT 0.210 1.078 0.851 1.280 ;
      RECT 0.000 1.120 0.210 1.280 ;
     END
  END VDD
END NAND2X2

MACRO MXI4X2
  CLASS CORE ;
  FOREIGN MXI4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.087 0.183 4.148 1.007 ;
      RECT 4.052 0.183 4.087 0.376 ;
      RECT 4.082 0.627 4.087 1.007 ;
      RECT 4.049 0.665 4.082 1.007 ;
      RECT 3.887 0.665 4.049 0.767 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.187 0.433 3.371 0.524 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.053 0.433 1.188 0.567 ;
     END
  END S0

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.437 0.302 1.548 0.533 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.292 0.300 2.413 0.367 ;
      RECT 2.233 0.300 2.292 0.561 ;
      RECT 2.231 0.306 2.233 0.561 ;
      RECT 2.205 0.474 2.231 0.561 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.969 0.306 0.993 0.361 ;
      RECT 0.908 0.306 0.969 0.527 ;
      RECT 0.862 0.450 0.908 0.527 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.526 0.209 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.924 -0.080 4.200 0.080 ;
      RECT 3.834 -0.080 3.924 0.122 ;
      RECT 3.468 -0.080 3.834 0.080 ;
      RECT 3.378 -0.080 3.468 0.122 ;
      RECT 2.360 -0.080 3.378 0.080 ;
      RECT 2.270 -0.080 2.360 0.217 ;
      RECT 1.522 -0.080 2.270 0.080 ;
      RECT 1.432 -0.080 1.522 0.217 ;
      RECT 1.042 -0.080 1.432 0.080 ;
      RECT 0.952 -0.080 1.042 0.220 ;
      RECT 0.151 -0.080 0.952 0.080 ;
      RECT 0.061 -0.080 0.151 0.329 ;
      RECT 0.000 -0.080 0.061 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.900 1.120 4.200 1.280 ;
      RECT 3.810 1.078 3.900 1.280 ;
      RECT 3.434 1.120 3.810 1.280 ;
      RECT 3.344 1.078 3.434 1.280 ;
      RECT 2.360 1.120 3.344 1.280 ;
      RECT 2.270 1.078 2.360 1.280 ;
      RECT 1.469 1.120 2.270 1.280 ;
      RECT 1.379 0.954 1.469 1.280 ;
      RECT 1.042 1.120 1.379 1.280 ;
      RECT 0.952 0.954 1.042 1.280 ;
      RECT 0.151 1.120 0.952 1.280 ;
      RECT 0.061 0.745 0.151 1.280 ;
      RECT 0.000 1.120 0.061 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.975 0.496 4.004 0.577 ;
      RECT 3.914 0.198 3.975 0.577 ;
      RECT 3.310 0.198 3.914 0.252 ;
      RECT 3.716 0.542 3.777 1.008 ;
      RECT 3.509 0.313 3.717 0.368 ;
      RECT 3.680 0.542 3.716 0.596 ;
      RECT 1.645 0.954 3.716 1.008 ;
      RECT 3.605 0.514 3.680 0.596 ;
      RECT 3.509 0.761 3.639 0.854 ;
      RECT 3.590 0.514 3.605 0.595 ;
      RECT 3.448 0.313 3.509 0.854 ;
      RECT 2.986 0.799 3.448 0.854 ;
      RECT 3.249 0.163 3.310 0.252 ;
      RECT 3.177 0.637 3.273 0.735 ;
      RECT 2.768 0.163 3.249 0.218 ;
      RECT 3.106 0.637 3.177 0.692 ;
      RECT 3.106 0.313 3.166 0.368 ;
      RECT 3.045 0.313 3.106 0.692 ;
      RECT 3.011 0.445 3.045 0.545 ;
      RECT 2.934 0.767 2.986 0.854 ;
      RECT 2.934 0.287 2.955 0.374 ;
      RECT 2.873 0.287 2.934 0.854 ;
      RECT 2.754 0.796 2.780 0.877 ;
      RECT 2.754 0.163 2.768 0.343 ;
      RECT 2.707 0.163 2.754 0.877 ;
      RECT 2.693 0.262 2.707 0.877 ;
      RECT 2.678 0.262 2.693 0.343 ;
      RECT 2.528 0.177 2.589 0.877 ;
      RECT 2.477 0.177 2.528 0.232 ;
      RECT 2.401 0.495 2.462 0.898 ;
      RECT 1.990 0.843 2.401 0.898 ;
      RECT 2.067 0.252 2.128 0.776 ;
      RECT 1.929 0.252 1.990 0.898 ;
      RECT 1.851 0.252 1.929 0.333 ;
      RECT 1.787 0.843 1.929 0.898 ;
      RECT 1.791 0.436 1.852 0.774 ;
      RECT 1.739 0.436 1.791 0.490 ;
      RECT 1.586 0.719 1.791 0.774 ;
      RECT 1.678 0.252 1.739 0.490 ;
      RECT 1.653 0.546 1.714 0.664 ;
      RECT 1.649 0.252 1.678 0.333 ;
      RECT 1.330 0.610 1.653 0.664 ;
      RECT 1.584 0.830 1.645 1.008 ;
      RECT 0.481 0.830 1.584 0.885 ;
      RECT 1.269 0.287 1.330 0.744 ;
      RECT 1.169 0.287 1.269 0.342 ;
      RECT 0.927 0.689 1.269 0.744 ;
      RECT 0.866 0.595 0.927 0.744 ;
      RECT 0.757 0.595 0.866 0.650 ;
      RECT 0.772 0.260 0.801 0.340 ;
      RECT 0.619 0.705 0.782 0.760 ;
      RECT 0.711 0.260 0.772 0.439 ;
      RECT 0.696 0.510 0.757 0.650 ;
      RECT 0.619 0.385 0.711 0.439 ;
      RECT 0.558 0.385 0.619 0.760 ;
      RECT 0.481 0.237 0.570 0.318 ;
      RECT 0.420 0.237 0.481 0.885 ;
      RECT 0.282 0.263 0.343 0.817 ;
  END
END MXI4X2

MACRO MXI2X2
  CLASS CORE ;
  FOREIGN MXI2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.400 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.883 0.293 0.944 0.888 ;
      RECT 0.838 0.833 0.883 0.888 ;
      RECT 0.716 0.833 0.838 1.005 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.179 0.656 0.313 0.767 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.387 0.506 0.493 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.252 0.433 1.363 0.576 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.352 -0.080 1.400 0.080 ;
      RECT 1.262 -0.080 1.352 0.122 ;
      RECT 0.459 -0.080 1.262 0.080 ;
      RECT 0.369 -0.080 0.459 0.261 ;
      RECT 0.000 -0.080 0.369 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.352 1.120 1.400 1.280 ;
      RECT 1.262 0.757 1.352 1.280 ;
      RECT 0.377 1.120 1.262 1.280 ;
      RECT 0.286 0.853 0.377 1.280 ;
      RECT 0.000 1.120 0.286 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.128 0.336 1.189 0.790 ;
      RECT 1.115 0.736 1.128 0.790 ;
      RECT 1.025 0.736 1.115 0.960 ;
      RECT 1.005 0.163 1.066 0.571 ;
      RECT 0.615 0.163 1.005 0.218 ;
      RECT 0.761 0.326 0.822 0.763 ;
      RECT 0.677 0.326 0.761 0.407 ;
      RECT 0.583 0.708 0.761 0.763 ;
      RECT 0.615 0.517 0.696 0.607 ;
      RECT 0.554 0.163 0.615 0.607 ;
      RECT 0.493 0.708 0.583 1.013 ;
      RECT 0.257 0.387 0.554 0.442 ;
      RECT 0.196 0.257 0.257 0.442 ;
      RECT 0.167 0.257 0.196 0.348 ;
      RECT 0.109 0.293 0.167 0.348 ;
      RECT 0.109 0.836 0.138 0.917 ;
      RECT 0.048 0.293 0.109 0.917 ;
  END
END MXI2X2

MACRO MX2X2
  CLASS CORE ;
  FOREIGN MX2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.494 0.194 1.556 0.977 ;
      RECT 1.480 0.194 1.494 0.439 ;
      RECT 1.446 0.700 1.494 0.977 ;
      RECT 1.461 0.194 1.480 0.395 ;
     END
  END Y

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.302 0.706 0.475 0.761 ;
      RECT 0.225 0.706 0.302 0.795 ;
      RECT 0.210 0.714 0.225 0.795 ;
     END
  END S0

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.215 0.526 0.387 0.633 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.285 0.306 1.364 0.361 ;
      RECT 1.222 0.306 1.285 0.367 ;
      RECT 1.160 0.306 1.222 0.575 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 -0.080 1.600 0.080 ;
      RECT 1.244 -0.080 1.336 0.223 ;
      RECT 0.407 -0.080 1.244 0.080 ;
      RECT 0.315 -0.080 0.407 0.296 ;
      RECT 0.000 -0.080 0.315 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.323 1.120 1.600 1.280 ;
      RECT 1.231 1.078 1.323 1.280 ;
      RECT 0.407 1.120 1.231 1.280 ;
      RECT 0.315 0.890 0.407 1.280 ;
      RECT 0.000 1.120 0.315 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.385 0.485 1.415 0.595 ;
      RECT 1.323 0.485 1.385 0.994 ;
      RECT 0.941 0.939 1.323 0.994 ;
      RECT 1.020 0.279 1.081 0.858 ;
      RECT 0.879 0.267 0.941 0.994 ;
      RECT 0.843 0.267 0.879 0.321 ;
      RECT 0.770 0.836 0.879 0.917 ;
      RECT 0.752 0.240 0.843 0.321 ;
      RECT 0.739 0.396 0.801 0.761 ;
      RECT 0.667 0.396 0.739 0.451 ;
      RECT 0.642 0.706 0.739 0.761 ;
      RECT 0.605 0.190 0.667 0.451 ;
      RECT 0.599 0.520 0.661 0.606 ;
      RECT 0.580 0.706 0.642 0.915 ;
      RECT 0.547 0.190 0.605 0.245 ;
      RECT 0.527 0.520 0.599 0.575 ;
      RECT 0.465 0.370 0.527 0.575 ;
      RECT 0.140 0.370 0.465 0.425 ;
      RECT 0.125 0.858 0.145 0.939 ;
      RECT 0.125 0.348 0.140 0.429 ;
      RECT 0.063 0.348 0.125 0.939 ;
      RECT 0.048 0.348 0.063 0.429 ;
      RECT 0.054 0.858 0.063 0.939 ;

      LAYER Metal2 ;
      RECT 0.100 0.325 1.063 0.375 ;
      RECT 0.580 0.825 1.200 0.875 ;
  END
END MX2X2

MACRO INVX3
  CLASS CORE ;
  FOREIGN INVX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.399 0.295 0.489 0.913 ;
      RECT 0.139 0.295 0.399 0.376 ;
      RECT 0.387 0.700 0.399 0.900 ;
      RECT 0.139 0.773 0.387 0.854 ;
      RECT 0.049 0.215 0.139 0.408 ;
      RECT 0.049 0.720 0.139 0.913 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.493 0.266 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.341 -0.080 0.700 0.080 ;
      RECT 0.251 -0.080 0.341 0.122 ;
      RECT 0.000 -0.080 0.251 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.341 1.120 0.700 1.280 ;
      RECT 0.251 1.078 0.341 1.280 ;
      RECT 0.000 1.120 0.251 1.280 ;
     END
  END VDD
END INVX3

MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.488 0.183 0.558 0.715 ;
      RECT 0.442 0.183 0.488 0.376 ;
      RECT 0.465 0.627 0.488 0.715 ;
      RECT 0.327 0.661 0.465 0.715 ;
      RECT 0.224 0.661 0.327 0.854 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.150 0.433 0.395 0.574 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.267 -0.080 0.600 0.080 ;
      RECT 0.164 -0.080 0.267 0.361 ;
      RECT 0.000 -0.080 0.164 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.497 1.120 0.600 1.280 ;
      RECT 0.495 1.078 0.497 1.280 ;
      RECT 0.395 1.064 0.495 1.280 ;
      RECT 0.394 1.078 0.395 1.280 ;
      RECT 0.000 1.120 0.394 1.280 ;
     END
  END VDD
END INVX2

MACRO DFFX2
  CLASS CORE ;
  FOREIGN DFFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN QN
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.405 0.323 3.466 0.793 ;
      RECT 3.385 0.323 3.405 0.439 ;
      RECT 3.390 0.738 3.405 0.793 ;
      RECT 3.300 0.738 3.390 0.819 ;
      RECT 3.358 0.323 3.385 0.404 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.071 0.167 3.086 0.248 ;
      RECT 2.995 0.167 3.071 0.257 ;
      RECT 2.900 0.202 2.995 0.257 ;
      RECT 2.958 0.683 2.979 0.764 ;
      RECT 2.900 0.567 2.958 0.764 ;
      RECT 2.888 0.202 2.900 0.764 ;
      RECT 2.856 0.202 2.888 0.633 ;
      RECT 2.839 0.202 2.856 0.621 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.390 0.335 0.487 0.494 ;
      RECT 0.354 0.335 0.390 0.415 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 0.214 0.505 0.315 0.633 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.599 -0.080 3.700 0.080 ;
      RECT 3.508 -0.080 3.599 0.122 ;
      RECT 3.300 -0.080 3.508 0.080 ;
      RECT 3.209 -0.080 3.300 0.122 ;
      RECT 2.872 -0.080 3.209 0.080 ;
      RECT 2.782 -0.080 2.872 0.122 ;
      RECT 2.349 -0.080 2.782 0.080 ;
      RECT 2.258 -0.080 2.349 0.287 ;
      RECT 1.651 -0.080 2.258 0.080 ;
      RECT 1.560 -0.080 1.651 0.329 ;
      RECT 1.073 -0.080 1.560 0.080 ;
      RECT 0.982 -0.080 1.073 0.287 ;
      RECT 0.294 -0.080 0.982 0.080 ;
      RECT 0.203 -0.080 0.294 0.122 ;
      RECT 0.000 -0.080 0.203 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.540 1.120 3.700 1.280 ;
      RECT 3.449 1.078 3.540 1.280 ;
      RECT 3.182 1.120 3.449 1.280 ;
      RECT 3.091 1.078 3.182 1.280 ;
      RECT 2.654 1.120 3.091 1.280 ;
      RECT 2.186 1.078 2.654 1.280 ;
      RECT 1.572 1.120 2.186 1.280 ;
      RECT 1.482 1.078 1.572 1.280 ;
      RECT 1.209 1.120 1.482 1.280 ;
      RECT 1.119 1.078 1.209 1.280 ;
      RECT 0.387 1.120 1.119 1.280 ;
      RECT 0.296 1.065 0.387 1.280 ;
      RECT 0.000 1.120 0.296 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.320 0.957 3.334 1.038 ;
      RECT 3.244 0.951 3.320 1.038 ;
      RECT 3.237 0.951 3.244 1.006 ;
      RECT 3.175 0.368 3.237 1.006 ;
      RECT 2.995 0.368 3.175 0.423 ;
      RECT 2.979 0.951 3.175 1.006 ;
      RECT 3.053 0.544 3.114 0.874 ;
      RECT 2.663 0.819 3.053 0.874 ;
      RECT 2.950 0.951 2.979 1.040 ;
      RECT 2.888 0.929 2.950 1.040 ;
      RECT 2.573 0.929 2.888 0.983 ;
      RECT 2.601 0.423 2.663 0.874 ;
      RECT 2.563 0.423 2.601 0.477 ;
      RECT 2.411 0.800 2.601 0.874 ;
      RECT 2.501 0.275 2.563 0.477 ;
      RECT 2.432 0.560 2.523 0.640 ;
      RECT 2.472 0.275 2.501 0.427 ;
      RECT 2.170 0.373 2.472 0.427 ;
      RECT 2.188 0.573 2.432 0.627 ;
      RECT 2.381 0.800 2.411 0.881 ;
      RECT 2.320 0.800 2.381 0.943 ;
      RECT 1.910 0.888 2.320 0.943 ;
      RECT 2.126 0.573 2.188 0.752 ;
      RECT 2.109 0.276 2.170 0.427 ;
      RECT 1.949 0.698 2.126 0.752 ;
      RECT 2.008 0.276 2.109 0.331 ;
      RECT 1.917 0.250 2.008 0.331 ;
      RECT 1.925 0.671 1.949 0.752 ;
      RECT 1.863 0.425 1.925 0.752 ;
      RECT 1.849 0.819 1.910 1.018 ;
      RECT 1.476 0.425 1.863 0.480 ;
      RECT 1.858 0.671 1.863 0.752 ;
      RECT 1.690 0.698 1.858 0.752 ;
      RECT 1.564 0.535 1.765 0.589 ;
      RECT 1.628 0.698 1.690 1.008 ;
      RECT 0.960 0.954 1.628 1.008 ;
      RECT 1.503 0.535 1.564 0.899 ;
      RECT 1.253 0.844 1.503 0.899 ;
      RECT 1.414 0.263 1.454 0.344 ;
      RECT 1.414 0.625 1.423 0.706 ;
      RECT 1.352 0.150 1.414 0.706 ;
      RECT 1.317 0.150 1.352 0.205 ;
      RECT 1.332 0.625 1.352 0.706 ;
      RECT 1.251 0.540 1.253 0.899 ;
      RECT 1.192 0.226 1.251 0.899 ;
      RECT 1.189 0.226 1.192 0.598 ;
      RECT 0.957 0.517 1.189 0.598 ;
      RECT 0.896 0.370 1.116 0.425 ;
      RECT 0.898 0.926 0.960 1.008 ;
      RECT 0.884 0.926 0.898 1.006 ;
      RECT 0.834 0.368 0.896 0.857 ;
      RECT 0.881 0.926 0.884 0.988 ;
      RECT 0.773 0.926 0.881 0.981 ;
      RECT 0.793 0.368 0.834 0.425 ;
      RECT 0.731 0.219 0.793 0.425 ;
      RECT 0.711 0.671 0.773 0.981 ;
      RECT 0.710 0.219 0.731 0.274 ;
      RECT 0.634 0.671 0.711 0.726 ;
      RECT 0.529 0.926 0.711 0.981 ;
      RECT 0.619 0.193 0.710 0.274 ;
      RECT 0.634 0.329 0.649 0.410 ;
      RECT 0.573 0.329 0.634 0.726 ;
      RECT 0.558 0.329 0.573 0.410 ;
      RECT 0.467 0.858 0.529 0.981 ;
      RECT 0.350 0.858 0.467 0.913 ;
      RECT 0.243 0.719 0.350 0.913 ;
      RECT 0.152 0.733 0.243 0.788 ;
      RECT 0.091 0.319 0.152 0.788 ;
      RECT 0.048 0.319 0.091 0.400 ;
  END
END DFFX2

MACRO BUFX3
  CLASS CORE ;
  FOREIGN BUFX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.469 0.287 0.498 0.368 ;
      RECT 0.469 0.433 0.488 0.752 ;
      RECT 0.408 0.287 0.469 0.752 ;
      RECT 0.398 0.433 0.408 0.752 ;
      RECT 0.387 0.433 0.398 0.633 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.433 0.147 0.562 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.647 -0.080 0.700 0.080 ;
      RECT 0.557 -0.080 0.647 0.122 ;
      RECT 0.000 -0.080 0.557 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.286 1.120 0.700 1.280 ;
      RECT 0.196 1.078 0.286 1.280 ;
      RECT 0.000 1.120 0.196 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.296 0.470 0.325 0.551 ;
      RECT 0.235 0.270 0.296 0.751 ;
      RECT 0.138 0.270 0.235 0.325 ;
      RECT 0.138 0.696 0.235 0.751 ;
      RECT 0.048 0.244 0.138 0.325 ;
      RECT 0.048 0.696 0.138 0.777 ;
  END
END BUFX3

MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.623 0.439 0.643 0.494 ;
      RECT 0.562 0.357 0.623 0.710 ;
      RECT 0.525 0.357 0.562 0.412 ;
      RECT 0.514 0.655 0.562 0.710 ;
      RECT 0.435 0.331 0.525 0.412 ;
      RECT 0.424 0.655 0.514 0.736 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.037 0.418 0.236 0.538 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.323 -0.080 0.700 0.080 ;
      RECT 0.233 -0.080 0.323 0.122 ;
      RECT 0.000 -0.080 0.233 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 1.120 0.700 1.280 ;
      RECT 0.298 1.078 0.313 1.280 ;
      RECT 0.237 1.065 0.298 1.280 ;
      RECT 0.223 1.078 0.237 1.280 ;
      RECT 0.000 1.120 0.223 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.363 0.490 0.430 0.571 ;
      RECT 0.302 0.301 0.363 0.712 ;
      RECT 0.164 0.301 0.302 0.356 ;
      RECT 0.164 0.657 0.302 0.712 ;
      RECT 0.074 0.275 0.164 0.356 ;
      RECT 0.074 0.657 0.164 0.738 ;
  END
END BUFX2

MACRO AOI33X2
  CLASS CORE ;
  FOREIGN AOI33X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.181 0.192 2.242 0.787 ;
      RECT 2.161 0.192 2.181 0.306 ;
      RECT 1.272 0.732 2.181 0.787 ;
      RECT 0.946 0.192 2.161 0.246 ;
      RECT 0.885 0.192 0.946 0.352 ;
      RECT 0.541 0.298 0.885 0.352 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.969 0.679 1.071 0.760 ;
      RECT 0.188 0.705 0.969 0.760 ;
      RECT 0.126 0.573 0.188 0.760 ;
      RECT 0.058 0.573 0.126 0.627 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.827 0.595 0.878 0.650 ;
      RECT 0.765 0.439 0.827 0.650 ;
      RECT 0.294 0.595 0.765 0.650 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.477 0.439 0.578 0.540 ;
      RECT 0.411 0.439 0.477 0.494 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.037 0.301 2.099 0.481 ;
      RECT 1.198 0.301 2.037 0.356 ;
      RECT 1.137 0.301 1.198 0.554 ;
      RECT 1.119 0.439 1.137 0.494 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.815 0.411 1.876 0.574 ;
      RECT 1.413 0.411 1.815 0.465 ;
      RECT 1.351 0.411 1.413 0.640 ;
      RECT 1.296 0.573 1.351 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 0.525 1.732 0.633 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.146 -0.080 2.300 0.080 ;
      RECT 2.055 -0.080 2.146 0.122 ;
      RECT 1.138 -0.080 2.055 0.080 ;
      RECT 1.047 -0.080 1.138 0.122 ;
      RECT 0.139 -0.080 1.047 0.080 ;
      RECT 0.048 -0.080 0.139 0.403 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.997 1.120 2.300 1.280 ;
      RECT 0.906 0.984 0.997 1.280 ;
      RECT 0.654 1.120 0.906 1.280 ;
      RECT 0.563 0.984 0.654 1.280 ;
      RECT 0.311 1.120 0.563 1.280 ;
      RECT 0.220 0.984 0.311 1.280 ;
      RECT 0.000 1.120 0.220 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.132 0.896 2.224 0.977 ;
      RECT 1.878 0.910 2.132 0.964 ;
      RECT 1.787 0.896 1.878 0.977 ;
      RECT 1.535 0.910 1.787 0.964 ;
      RECT 1.444 0.896 1.535 0.977 ;
      RECT 1.192 0.910 1.444 0.964 ;
      RECT 1.162 0.896 1.192 0.977 ;
      RECT 1.100 0.814 1.162 0.977 ;
      RECT 0.048 0.814 1.100 0.869 ;
  END
END AOI33X2

MACRO AOI32X2
  CLASS CORE ;
  FOREIGN AOI32X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.877 0.348 1.941 0.789 ;
      RECT 1.857 0.348 1.877 0.439 ;
      RECT 1.756 0.735 1.877 0.789 ;
      RECT 1.727 0.348 1.857 0.402 ;
      RECT 1.663 0.721 1.756 0.802 ;
      RECT 1.664 0.281 1.727 0.402 ;
      RECT 0.894 0.281 1.664 0.336 ;
      RECT 1.404 0.732 1.663 0.787 ;
      RECT 1.310 0.719 1.404 0.800 ;
      RECT 0.831 0.189 0.894 0.336 ;
      RECT 0.556 0.189 0.831 0.244 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.241 0.606 1.742 0.661 ;
      RECT 1.178 0.439 1.241 0.661 ;
      RECT 1.150 0.439 1.178 0.507 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.466 0.433 1.598 0.507 ;
      RECT 1.372 0.433 1.466 0.550 ;
      RECT 1.371 0.433 1.372 0.507 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.993 0.569 1.056 0.692 ;
      RECT 0.948 0.626 0.993 0.692 ;
      RECT 0.178 0.637 0.948 0.692 ;
      RECT 0.114 0.573 0.178 0.692 ;
      RECT 0.059 0.573 0.114 0.627 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.766 0.439 0.872 0.577 ;
      RECT 0.302 0.523 0.766 0.577 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.554 0.413 0.584 0.468 ;
      RECT 0.490 0.306 0.554 0.468 ;
      RECT 0.423 0.306 0.490 0.361 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.884 -0.080 2.000 0.080 ;
      RECT 1.791 -0.080 1.884 0.275 ;
      RECT 1.168 -0.080 1.791 0.080 ;
      RECT 1.074 -0.080 1.168 0.122 ;
      RECT 0.128 -0.080 1.074 0.080 ;
      RECT 0.065 -0.080 0.128 0.325 ;
      RECT 0.000 -0.080 0.065 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.026 1.120 2.000 1.280 ;
      RECT 0.933 0.989 1.026 1.280 ;
      RECT 0.674 1.120 0.933 1.280 ;
      RECT 0.580 0.989 0.674 1.280 ;
      RECT 0.320 1.120 0.580 1.280 ;
      RECT 0.226 0.989 0.320 1.280 ;
      RECT 0.000 1.120 0.226 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.839 0.896 1.933 0.977 ;
      RECT 1.580 0.910 1.839 0.964 ;
      RECT 1.486 0.896 1.580 0.977 ;
      RECT 1.227 0.910 1.486 0.964 ;
      RECT 1.197 0.896 1.227 0.977 ;
      RECT 1.134 0.812 1.197 0.977 ;
      RECT 0.850 0.812 1.134 0.867 ;
      RECT 0.756 0.799 0.850 0.880 ;
      RECT 0.497 0.810 0.756 0.864 ;
      RECT 0.404 0.796 0.497 0.877 ;
      RECT 0.143 0.810 0.404 0.864 ;
      RECT 0.050 0.796 0.143 0.877 ;
  END
END AOI32X2

MACRO AOI31X2
  CLASS CORE ;
  FOREIGN AOI31X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.292 0.627 1.354 0.800 ;
      RECT 1.282 0.627 1.292 0.706 ;
      RECT 1.187 0.627 1.282 0.682 ;
      RECT 1.125 0.268 1.187 0.682 ;
      RECT 0.482 0.268 1.125 0.323 ;
      RECT 0.420 0.158 0.482 0.323 ;
      RECT 0.048 0.158 0.420 0.213 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.248 0.433 1.395 0.557 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.318 0.413 0.614 0.468 ;
      RECT 0.236 0.306 0.318 0.468 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.851 0.527 0.882 0.582 ;
      RECT 0.749 0.439 0.851 0.582 ;
      RECT 0.329 0.527 0.749 0.582 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.990 0.490 1.052 0.692 ;
      RECT 0.140 0.637 0.990 0.692 ;
      RECT 0.038 0.550 0.140 0.692 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.336 -0.080 1.600 0.080 ;
      RECT 1.331 -0.080 1.336 0.122 ;
      RECT 1.269 -0.080 1.331 0.304 ;
      RECT 1.244 -0.080 1.269 0.122 ;
      RECT 0.636 -0.080 1.244 0.080 ;
      RECT 0.544 -0.080 0.636 0.198 ;
      RECT 0.000 -0.080 0.544 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.002 1.120 1.600 1.280 ;
      RECT 0.910 0.911 1.002 1.280 ;
      RECT 0.657 1.120 0.910 1.280 ;
      RECT 0.566 0.911 0.657 1.280 ;
      RECT 0.312 1.120 0.566 1.280 ;
      RECT 0.221 0.911 0.312 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.129 0.910 1.541 0.964 ;
      RECT 1.067 0.746 1.129 0.964 ;
      RECT 0.048 0.746 1.067 0.801 ;
  END
END AOI31X2

MACRO AOI2BB2X2
  CLASS CORE ;
  FOREIGN AOI2BB2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.508 0.306 1.542 0.361 ;
      RECT 1.446 0.192 1.508 0.977 ;
      RECT 0.773 0.192 1.446 0.246 ;
      RECT 1.304 0.923 1.446 0.977 ;
      RECT 1.203 0.923 1.304 1.040 ;
      RECT 1.187 0.967 1.203 1.040 ;
      RECT 1.094 0.986 1.187 1.040 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.104 0.543 1.201 0.737 ;
      RECT 0.512 0.682 1.104 0.737 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.294 0.379 1.371 0.498 ;
      RECT 0.672 0.379 1.294 0.433 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.343 0.388 0.496 0.500 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.038 0.445 0.140 0.633 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.072 -0.080 1.600 0.080 ;
      RECT 0.980 -0.080 1.072 0.122 ;
      RECT 0.516 -0.080 0.980 0.080 ;
      RECT 0.424 -0.080 0.516 0.289 ;
      RECT 0.140 -0.080 0.424 0.080 ;
      RECT 0.048 -0.080 0.140 0.122 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.541 1.120 1.600 1.280 ;
      RECT 1.449 1.078 1.541 1.280 ;
      RECT 0.840 1.120 1.449 1.280 ;
      RECT 0.749 0.988 0.840 1.280 ;
      RECT 0.496 1.120 0.749 1.280 ;
      RECT 0.404 0.988 0.496 1.280 ;
      RECT 0.000 1.120 0.404 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.576 0.808 1.358 0.863 ;
      RECT 0.276 0.571 0.991 0.626 ;
      RECT 0.214 0.288 0.276 0.788 ;
      RECT 0.048 0.733 0.214 0.788 ;
  END
END AOI2BB2X2

MACRO AOI2BB1X2
  CLASS CORE ;
  FOREIGN AOI2BB1X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.147 0.323 1.211 0.765 ;
      RECT 0.803 0.323 1.147 0.377 ;
      RECT 0.868 0.711 1.147 0.765 ;
      RECT 0.833 0.711 0.868 0.894 ;
      RECT 0.737 0.711 0.833 0.904 ;
      RECT 0.739 0.300 0.803 0.377 ;
      RECT 0.674 0.162 0.739 0.377 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.009 0.439 1.073 0.638 ;
      RECT 0.671 0.439 1.009 0.494 ;
      RECT 0.606 0.439 0.671 0.538 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.194 0.555 0.387 0.652 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.300 0.149 0.429 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.968 -0.080 1.300 0.080 ;
      RECT 0.872 -0.080 0.968 0.122 ;
      RECT 0.552 -0.080 0.872 0.080 ;
      RECT 0.456 -0.080 0.552 0.198 ;
      RECT 0.146 -0.080 0.456 0.080 ;
      RECT 0.051 -0.080 0.146 0.198 ;
      RECT 0.000 -0.080 0.051 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.193 1.120 1.300 1.280 ;
      RECT 1.097 0.860 1.193 1.280 ;
      RECT 0.461 1.120 1.097 1.280 ;
      RECT 0.366 1.078 0.461 1.280 ;
      RECT 0.000 1.120 0.366 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.518 0.596 0.900 0.651 ;
      RECT 0.453 0.427 0.518 0.762 ;
      RECT 0.333 0.427 0.453 0.482 ;
      RECT 0.146 0.707 0.453 0.762 ;
      RECT 0.269 0.183 0.333 0.482 ;
      RECT 0.051 0.707 0.146 0.900 ;
  END
END AOI2BB1X2

MACRO AOI22X2
  CLASS CORE ;
  FOREIGN AOI22X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.480 0.321 1.542 0.761 ;
      RECT 0.393 0.321 1.480 0.376 ;
      RECT 1.368 0.706 1.480 0.761 ;
      RECT 1.302 0.706 1.368 0.789 ;
      RECT 0.932 0.735 1.302 0.789 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.653 0.456 0.715 0.575 ;
      RECT 0.298 0.456 0.653 0.511 ;
      RECT 0.246 0.439 0.298 0.511 ;
      RECT 0.185 0.439 0.246 0.562 ;
      RECT 0.113 0.493 0.185 0.562 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.329 0.573 0.475 0.663 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.356 0.438 1.418 0.551 ;
      RECT 1.009 0.438 1.356 0.493 ;
      RECT 0.944 0.438 1.009 0.494 ;
      RECT 0.882 0.438 0.944 0.664 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.061 0.567 1.207 0.661 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.444 -0.080 1.600 0.080 ;
      RECT 1.352 -0.080 1.444 0.122 ;
      RECT 0.787 -0.080 1.352 0.080 ;
      RECT 0.695 -0.080 0.787 0.122 ;
      RECT 0.140 -0.080 0.695 0.080 ;
      RECT 0.048 -0.080 0.140 0.305 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.657 1.120 1.600 1.280 ;
      RECT 0.566 0.888 0.657 1.280 ;
      RECT 0.312 1.120 0.566 1.280 ;
      RECT 0.221 0.888 0.312 1.280 ;
      RECT 0.000 1.120 0.221 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.815 0.886 1.541 0.940 ;
      RECT 0.815 0.732 0.830 0.787 ;
      RECT 0.753 0.732 0.815 0.940 ;
      RECT 0.048 0.732 0.753 0.787 ;
  END
END AOI22X2

MACRO AOI222X2
  CLASS CORE ;
  FOREIGN AOI222X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.500 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.336 0.268 2.399 0.743 ;
      RECT 2.263 0.268 2.336 0.367 ;
      RECT 2.263 0.688 2.336 0.743 ;
      RECT 2.024 0.268 2.263 0.323 ;
      RECT 2.201 0.688 2.263 0.761 ;
      RECT 1.797 0.688 2.201 0.743 ;
      RECT 1.905 0.249 2.024 0.323 ;
      RECT 1.318 0.268 1.905 0.323 ;
      RECT 1.190 0.249 1.318 0.323 ;
      RECT 0.395 0.268 1.190 0.323 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.628 0.556 0.725 0.620 ;
      RECT 0.299 0.565 0.628 0.620 ;
      RECT 0.156 0.565 0.299 0.627 ;
      RECT 0.093 0.521 0.156 0.627 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.319 0.398 0.517 0.507 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.951 0.439 1.558 0.494 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.130 0.558 1.331 0.627 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.210 0.439 2.273 0.545 ;
      RECT 1.665 0.439 2.210 0.494 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.814 0.556 2.016 0.627 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.353 -0.080 2.500 0.080 ;
      RECT 2.261 -0.080 2.353 0.198 ;
      RECT 1.659 -0.080 2.261 0.080 ;
      RECT 1.567 -0.080 1.659 0.198 ;
      RECT 0.874 -0.080 1.567 0.080 ;
      RECT 0.782 -0.080 0.874 0.198 ;
      RECT 0.141 -0.080 0.782 0.080 ;
      RECT 0.049 -0.080 0.141 0.275 ;
      RECT 0.000 -0.080 0.049 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.833 1.120 2.500 1.280 ;
      RECT 0.741 0.911 0.833 1.280 ;
      RECT 0.487 1.120 0.741 1.280 ;
      RECT 0.395 0.911 0.487 1.280 ;
      RECT 0.141 1.120 0.395 1.280 ;
      RECT 0.049 0.911 0.141 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.931 0.910 2.408 0.964 ;
      RECT 0.222 0.688 1.542 0.743 ;
  END
END AOI222X2

MACRO AOI221X2
  CLASS CORE ;
  FOREIGN AOI221X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.807 0.312 1.868 0.836 ;
      RECT 1.457 0.312 1.807 0.367 ;
      RECT 1.761 0.755 1.807 0.836 ;
      RECT 1.391 0.300 1.457 0.367 ;
      RECT 1.330 0.225 1.391 0.367 ;
      RECT 0.387 0.225 1.330 0.280 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.678 0.439 1.739 0.543 ;
      RECT 1.457 0.439 1.678 0.494 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.663 0.493 0.711 0.558 ;
      RECT 0.562 0.433 0.663 0.558 ;
      RECT 0.077 0.504 0.562 0.558 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.313 0.375 0.414 0.430 ;
      RECT 0.212 0.306 0.313 0.430 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.993 0.595 1.572 0.650 ;
      RECT 0.932 0.573 0.993 0.650 ;
      RECT 0.917 0.595 0.932 0.650 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.087 0.396 1.233 0.500 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.636 -0.080 2.100 0.080 ;
      RECT 1.546 -0.080 1.636 0.198 ;
      RECT 0.870 -0.080 1.546 0.080 ;
      RECT 0.780 -0.080 0.870 0.122 ;
      RECT 0.138 -0.080 0.780 0.080 ;
      RECT 0.048 -0.080 0.138 0.198 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.817 1.120 2.100 1.280 ;
      RECT 0.727 0.903 0.817 1.280 ;
      RECT 0.477 1.120 0.727 1.280 ;
      RECT 0.387 0.903 0.477 1.280 ;
      RECT 0.138 1.120 0.387 1.280 ;
      RECT 0.048 0.903 0.138 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.912 0.962 2.020 1.017 ;
      RECT 0.944 0.768 1.511 0.823 ;
      RECT 0.883 0.707 0.944 0.823 ;
      RECT 0.217 0.707 0.883 0.762 ;
  END
END AOI221X2

MACRO AOI21X2
  CLASS CORE ;
  FOREIGN AOI21X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.030 0.345 1.095 0.789 ;
      RECT 0.867 0.345 1.030 0.400 ;
      RECT 0.989 0.706 1.030 0.789 ;
      RECT 0.974 0.735 0.989 0.789 ;
      RECT 0.771 0.268 0.867 0.400 ;
      RECT 0.300 0.345 0.771 0.400 ;
      RECT 0.235 0.294 0.300 0.400 ;
      RECT 0.146 0.294 0.235 0.349 ;
      RECT 0.051 0.268 0.146 0.349 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.830 0.485 0.936 0.627 ;
      RECT 0.803 0.573 0.830 0.627 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.311 0.595 0.518 0.669 ;
      RECT 0.246 0.573 0.311 0.669 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.146 0.457 0.763 0.512 ;
      RECT 0.039 0.433 0.146 0.530 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.082 -0.080 1.300 0.080 ;
      RECT 0.986 -0.080 1.082 0.122 ;
      RECT 0.506 -0.080 0.986 0.080 ;
      RECT 0.411 -0.080 0.506 0.275 ;
      RECT 0.000 -0.080 0.411 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.687 1.120 1.300 1.280 ;
      RECT 0.591 0.888 0.687 1.280 ;
      RECT 0.326 1.120 0.591 1.280 ;
      RECT 0.231 0.888 0.326 1.280 ;
      RECT 0.000 1.120 0.231 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.154 0.873 1.249 0.954 ;
      RECT 0.871 0.873 1.154 0.927 ;
      RECT 0.806 0.732 0.871 0.927 ;
      RECT 0.051 0.732 0.806 0.787 ;
  END
END AOI21X2

MACRO AND4X2
  CLASS CORE ;
  FOREIGN AND4X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.100 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.049 0.700 1.061 0.767 ;
      RECT 1.031 0.358 1.049 0.767 ;
      RECT 0.985 0.199 1.031 0.964 ;
      RECT 0.967 0.199 0.985 0.413 ;
      RECT 0.967 0.648 0.985 0.964 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.694 0.524 0.733 0.606 ;
      RECT 0.610 0.439 0.694 0.606 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.478 0.581 0.542 0.761 ;
      RECT 0.426 0.706 0.478 0.761 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.279 0.537 0.358 0.646 ;
      RECT 0.222 0.537 0.279 0.645 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.039 0.398 0.157 0.556 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.815 -0.080 1.100 0.080 ;
      RECT 0.721 -0.080 0.815 0.122 ;
      RECT 0.000 -0.080 0.721 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.838 1.120 1.100 1.280 ;
      RECT 0.724 1.064 0.838 1.280 ;
      RECT 0.514 1.120 0.724 1.280 ;
      RECT 0.419 1.078 0.514 1.280 ;
      RECT 0.158 1.120 0.419 1.280 ;
      RECT 0.049 1.078 0.158 1.280 ;
      RECT 0.000 1.120 0.049 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.889 0.473 0.919 0.556 ;
      RECT 0.825 0.211 0.889 0.889 ;
      RECT 0.156 0.211 0.825 0.265 ;
      RECT 0.208 0.835 0.825 0.889 ;
      RECT 0.076 0.211 0.156 0.343 ;
      RECT 0.061 0.250 0.076 0.343 ;
  END
END AND4X2

MACRO AOI211X2
  CLASS CORE ;
  FOREIGN AOI211X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.600 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.471 0.249 1.533 0.761 ;
      RECT 1.414 0.249 1.471 0.304 ;
      RECT 1.177 0.706 1.471 0.761 ;
      RECT 1.323 0.223 1.414 0.304 ;
      RECT 0.980 0.236 1.323 0.290 ;
      RECT 1.100 0.706 1.177 0.807 ;
      RECT 1.086 0.726 1.100 0.807 ;
      RECT 0.762 0.223 0.980 0.304 ;
      RECT 0.749 0.223 0.762 0.290 ;
      RECT 0.143 0.236 0.749 0.290 ;
      RECT 0.051 0.223 0.143 0.304 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.345 0.365 1.407 0.539 ;
      RECT 1.282 0.365 1.345 0.439 ;
      RECT 0.905 0.365 1.282 0.420 ;
      RECT 0.843 0.365 0.905 0.627 ;
      RECT 0.769 0.550 0.843 0.627 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.021 0.550 1.207 0.645 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.236 0.539 0.399 0.627 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.601 0.494 0.615 0.621 ;
      RECT 0.539 0.399 0.601 0.621 ;
      RECT 0.207 0.399 0.539 0.454 ;
      RECT 0.524 0.540 0.539 0.621 ;
      RECT 0.120 0.386 0.207 0.467 ;
      RECT 0.116 0.386 0.120 0.494 ;
      RECT 0.058 0.399 0.116 0.494 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.208 -0.080 1.600 0.080 ;
      RECT 1.116 -0.080 1.208 0.122 ;
      RECT 0.498 -0.080 1.116 0.080 ;
      RECT 0.407 -0.080 0.498 0.122 ;
      RECT 0.000 -0.080 0.407 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.659 1.120 1.600 1.280 ;
      RECT 0.567 0.925 0.659 1.280 ;
      RECT 0.314 1.120 0.567 1.280 ;
      RECT 0.222 0.925 0.314 1.280 ;
      RECT 0.000 1.120 0.222 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.430 0.881 1.522 0.962 ;
      RECT 0.937 0.894 1.430 0.949 ;
      RECT 0.875 0.688 0.937 0.949 ;
      RECT 0.050 0.688 0.875 0.743 ;
  END
END AOI211X2

MACRO AND3X2
  CLASS CORE ;
  FOREIGN AND3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.807 0.317 0.845 0.761 ;
      RECT 0.783 0.188 0.807 0.761 ;
      RECT 0.715 0.188 0.783 0.383 ;
      RECT 0.768 0.652 0.783 0.761 ;
      RECT 0.753 0.652 0.768 0.733 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.510 0.600 0.540 0.689 ;
      RECT 0.447 0.433 0.510 0.689 ;
      RECT 0.398 0.433 0.447 0.500 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.280 0.564 0.342 0.689 ;
      RECT 0.218 0.567 0.280 0.689 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.142 0.587 0.155 0.668 ;
      RECT 0.038 0.587 0.142 0.773 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.600 -0.080 0.900 0.080 ;
      RECT 0.507 -0.080 0.600 0.122 ;
      RECT 0.000 -0.080 0.507 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.638 1.120 0.900 1.280 ;
      RECT 0.545 1.065 0.638 1.280 ;
      RECT 0.000 1.120 0.545 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.675 0.488 0.720 0.583 ;
      RECT 0.652 0.488 0.675 0.829 ;
      RECT 0.612 0.324 0.652 0.829 ;
      RECT 0.589 0.324 0.612 0.543 ;
      RECT 0.305 0.774 0.612 0.829 ;
      RECT 0.142 0.324 0.589 0.379 ;
      RECT 0.243 0.774 0.305 1.008 ;
      RECT 0.142 0.954 0.243 1.008 ;
      RECT 0.049 0.298 0.142 0.379 ;
      RECT 0.048 0.954 0.142 1.049 ;
  END
END AND3X2

MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.642 0.227 0.654 0.767 ;
      RECT 0.593 0.195 0.642 1.002 ;
      RECT 0.582 0.195 0.593 0.439 ;
      RECT 0.552 0.688 0.593 1.002 ;
      RECT 0.552 0.195 0.582 0.390 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.212 0.833 0.361 0.935 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.138 0.504 0.202 0.585 ;
      RECT 0.037 0.504 0.138 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.440 -0.080 0.700 0.080 ;
      RECT 0.350 -0.080 0.440 0.122 ;
      RECT 0.000 -0.080 0.350 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.151 1.120 0.700 1.280 ;
      RECT 0.048 1.078 0.151 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.325 0.512 0.521 0.594 ;
      RECT 0.264 0.348 0.325 0.737 ;
      RECT 0.138 0.348 0.264 0.402 ;
      RECT 0.216 0.654 0.264 0.737 ;
      RECT 0.048 0.321 0.138 0.402 ;
  END
END AND2X2

MACRO ADDHX2
  CLASS CORE ;
  FOREIGN ADDHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.200 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.539 0.306 1.601 0.392 ;
      RECT 1.142 0.674 1.578 0.755 ;
      RECT 0.947 0.319 1.539 0.374 ;
      RECT 1.009 0.687 1.142 0.755 ;
      RECT 0.879 0.687 1.009 0.761 ;
      RECT 0.894 0.306 0.947 0.374 ;
      RECT 0.879 0.306 0.894 0.387 ;
      RECT 0.818 0.306 0.879 0.761 ;
      RECT 0.803 0.306 0.818 0.387 ;
      RECT 0.812 0.669 0.818 0.761 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.985 0.324 3.099 0.405 ;
      RECT 2.964 0.324 2.985 0.439 ;
      RECT 2.967 0.626 2.982 0.733 ;
      RECT 2.964 0.626 2.967 0.761 ;
      RECT 2.902 0.350 2.964 0.761 ;
      RECT 2.890 0.626 2.902 0.733 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.386 0.438 1.477 0.519 ;
      RECT 1.364 0.438 1.386 0.506 ;
      RECT 1.302 0.439 1.364 0.506 ;
      RECT 1.104 0.451 1.302 0.506 ;
      RECT 1.042 0.451 1.104 0.619 ;
      RECT 1.013 0.538 1.042 0.619 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.253 0.454 2.525 0.535 ;
      RECT 2.191 0.439 2.253 0.535 ;
      RECT 2.054 0.454 2.191 0.535 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.905 -0.080 3.200 0.080 ;
      RECT 2.813 -0.080 2.905 0.211 ;
      RECT 2.566 -0.080 2.813 0.080 ;
      RECT 2.474 -0.080 2.566 0.220 ;
      RECT 2.221 -0.080 2.474 0.080 ;
      RECT 2.129 -0.080 2.221 0.220 ;
      RECT 0.496 -0.080 2.129 0.080 ;
      RECT 0.404 -0.080 0.496 0.122 ;
      RECT 0.140 -0.080 0.404 0.080 ;
      RECT 0.048 -0.080 0.140 0.215 ;
      RECT 0.000 -0.080 0.048 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.809 1.120 3.200 1.280 ;
      RECT 2.718 0.989 2.809 1.280 ;
      RECT 2.448 1.120 2.718 1.280 ;
      RECT 2.357 0.989 2.448 1.280 ;
      RECT 2.104 1.120 2.357 1.280 ;
      RECT 2.012 1.002 2.104 1.280 ;
      RECT 1.767 1.120 2.012 1.280 ;
      RECT 1.675 1.065 1.767 1.280 ;
      RECT 0.496 1.120 1.675 1.280 ;
      RECT 0.404 1.078 0.496 1.280 ;
      RECT 0.140 1.120 0.404 1.280 ;
      RECT 0.048 1.002 0.140 1.280 ;
      RECT 0.000 1.120 0.048 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.760 0.514 2.789 0.595 ;
      RECT 2.698 0.514 2.760 0.658 ;
      RECT 2.646 0.313 2.738 0.394 ;
      RECT 1.918 0.604 2.698 0.658 ;
      RECT 1.996 0.324 2.646 0.379 ;
      RECT 2.246 0.713 2.621 0.794 ;
      RECT 2.185 0.713 2.246 0.896 ;
      RECT 1.725 0.842 2.185 0.896 ;
      RECT 1.934 0.158 1.996 0.379 ;
      RECT 1.725 0.158 1.934 0.213 ;
      RECT 1.851 0.604 1.918 0.762 ;
      RECT 1.826 0.289 1.851 0.762 ;
      RECT 1.789 0.289 1.826 0.658 ;
      RECT 1.663 0.158 1.725 0.896 ;
      RECT 1.352 0.158 1.663 0.213 ;
      RECT 1.538 0.842 1.663 0.896 ;
      RECT 1.476 0.842 1.538 1.024 ;
      RECT 1.406 0.969 1.476 1.024 ;
      RECT 1.314 0.969 1.406 1.050 ;
      RECT 0.637 0.995 1.314 1.050 ;
      RECT 0.620 0.158 1.067 0.213 ;
      RECT 0.793 0.885 1.061 0.939 ;
      RECT 0.731 0.843 0.793 0.939 ;
      RECT 0.675 0.302 0.737 0.733 ;
      RECT 0.388 0.843 0.731 0.898 ;
      RECT 0.609 0.302 0.675 0.357 ;
      RECT 0.609 0.652 0.675 0.733 ;
      RECT 0.575 0.952 0.637 1.050 ;
      RECT 0.558 0.158 0.620 0.248 ;
      RECT 0.264 0.952 0.575 1.007 ;
      RECT 0.388 0.193 0.558 0.248 ;
      RECT 0.326 0.193 0.388 0.898 ;
      RECT 0.221 0.325 0.326 0.406 ;
      RECT 0.221 0.652 0.326 0.733 ;
      RECT 0.202 0.850 0.264 1.007 ;
      RECT 0.156 0.505 0.248 0.586 ;
      RECT 0.133 0.850 0.202 0.905 ;
      RECT 0.133 0.531 0.156 0.586 ;
      RECT 0.071 0.531 0.133 0.905 ;
  END
END ADDHX2

MACRO ADDFX2
  CLASS CORE ;
  FOREIGN ADDFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.700 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.557 0.306 3.569 0.424 ;
      RECT 3.557 0.665 3.565 0.746 ;
      RECT 3.496 0.306 3.557 0.746 ;
      RECT 3.478 0.306 3.496 0.424 ;
      RECT 3.474 0.665 3.496 0.746 ;
      RECT 3.405 0.306 3.478 0.361 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.139 0.340 3.205 0.421 ;
      RECT 3.139 0.665 3.199 0.746 ;
      RECT 3.078 0.340 3.139 0.746 ;
      RECT 3.053 0.573 3.078 0.627 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.461 0.433 2.532 0.488 ;
      RECT 2.400 0.433 2.461 0.767 ;
      RECT 2.296 0.682 2.400 0.767 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.119 0.486 0.203 0.567 ;
      RECT 0.112 0.486 0.119 0.627 ;
      RECT 0.057 0.512 0.112 0.627 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.040 0.560 1.291 0.640 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.388 -0.080 3.700 0.080 ;
      RECT 3.297 -0.080 3.388 0.122 ;
      RECT 2.691 -0.080 3.297 0.080 ;
      RECT 2.600 -0.080 2.691 0.122 ;
      RECT 1.261 -0.080 2.600 0.080 ;
      RECT 1.171 -0.080 1.261 0.199 ;
      RECT 0.343 -0.080 1.171 0.080 ;
      RECT 0.252 -0.080 0.343 0.122 ;
      RECT 0.000 -0.080 0.252 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.384 1.120 3.700 1.280 ;
      RECT 3.293 1.078 3.384 1.280 ;
      RECT 2.385 1.120 3.293 1.280 ;
      RECT 2.294 1.078 2.385 1.280 ;
      RECT 0.320 1.120 2.294 1.280 ;
      RECT 0.230 1.078 0.320 1.280 ;
      RECT 0.000 1.120 0.230 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.373 0.480 3.434 0.569 ;
      RECT 3.341 0.514 3.373 0.569 ;
      RECT 3.280 0.514 3.341 0.939 ;
      RECT 2.791 0.885 3.280 0.939 ;
      RECT 2.508 0.995 3.034 1.050 ;
      RECT 2.971 0.150 3.013 0.205 ;
      RECT 2.971 0.743 2.983 0.824 ;
      RECT 2.910 0.150 2.971 0.824 ;
      RECT 2.535 0.193 2.910 0.248 ;
      RECT 2.892 0.743 2.910 0.824 ;
      RECT 2.790 0.320 2.848 0.562 ;
      RECT 2.790 0.765 2.791 0.939 ;
      RECT 2.787 0.320 2.790 0.939 ;
      RECT 2.730 0.507 2.787 0.939 ;
      RECT 2.728 0.507 2.730 0.846 ;
      RECT 2.700 0.765 2.728 0.846 ;
      RECT 2.595 0.302 2.656 0.685 ;
      RECT 2.412 0.302 2.595 0.357 ;
      RECT 2.584 0.630 2.595 0.685 ;
      RECT 2.523 0.630 2.584 0.846 ;
      RECT 2.473 0.150 2.535 0.248 ;
      RECT 2.447 0.954 2.508 1.050 ;
      RECT 1.570 0.150 2.473 0.205 ;
      RECT 2.097 0.954 2.447 1.008 ;
      RECT 2.351 0.260 2.412 0.357 ;
      RECT 1.781 0.260 2.351 0.314 ;
      RECT 2.288 0.523 2.339 0.604 ;
      RECT 2.226 0.377 2.288 0.604 ;
      RECT 2.220 0.549 2.226 0.604 ;
      RECT 2.158 0.549 2.220 0.898 ;
      RECT 2.096 0.852 2.097 1.008 ;
      RECT 2.036 0.377 2.096 1.008 ;
      RECT 2.034 0.377 2.036 0.907 ;
      RECT 1.915 0.852 2.034 0.907 ;
      RECT 1.911 0.426 1.973 0.798 ;
      RECT 1.903 0.426 1.911 0.481 ;
      RECT 1.814 0.743 1.911 0.798 ;
      RECT 1.842 0.377 1.903 0.481 ;
      RECT 1.781 0.562 1.850 0.643 ;
      RECT 1.785 0.743 1.814 0.915 ;
      RECT 1.753 0.743 1.785 1.050 ;
      RECT 1.719 0.260 1.781 0.688 ;
      RECT 1.723 0.835 1.753 1.050 ;
      RECT 1.403 0.965 1.723 1.050 ;
      RECT 1.648 0.632 1.719 0.688 ;
      RECT 1.415 0.493 1.658 0.576 ;
      RECT 1.622 0.632 1.648 0.815 ;
      RECT 1.587 0.632 1.622 0.829 ;
      RECT 1.539 0.748 1.587 0.829 ;
      RECT 1.508 0.150 1.570 0.417 ;
      RECT 1.531 0.748 1.539 0.911 ;
      RECT 1.478 0.761 1.531 0.911 ;
      RECT 1.479 0.270 1.508 0.417 ;
      RECT 1.109 0.270 1.479 0.325 ;
      RECT 0.918 0.856 1.478 0.911 ;
      RECT 1.353 0.389 1.415 0.801 ;
      RECT 0.443 0.995 1.403 1.050 ;
      RECT 0.986 0.389 1.353 0.444 ;
      RECT 1.041 0.746 1.353 0.801 ;
      RECT 1.048 0.208 1.109 0.325 ;
      RECT 0.654 0.208 1.048 0.263 ;
      RECT 0.980 0.710 1.041 0.801 ;
      RECT 0.925 0.343 0.986 0.444 ;
      RECT 0.857 0.721 0.918 0.911 ;
      RECT 0.849 0.721 0.857 0.776 ;
      RECT 0.788 0.494 0.849 0.776 ;
      RECT 0.734 0.832 0.796 0.940 ;
      RECT 0.777 0.494 0.788 0.549 ;
      RECT 0.715 0.338 0.777 0.549 ;
      RECT 0.567 0.832 0.734 0.887 ;
      RECT 0.654 0.604 0.699 0.752 ;
      RECT 0.638 0.208 0.654 0.752 ;
      RECT 0.593 0.208 0.638 0.658 ;
      RECT 0.531 0.726 0.567 0.887 ;
      RECT 0.506 0.332 0.531 0.887 ;
      RECT 0.470 0.332 0.506 0.781 ;
      RECT 0.402 0.700 0.470 0.781 ;
      RECT 0.382 0.870 0.443 1.050 ;
      RECT 0.368 0.486 0.398 0.567 ;
      RECT 0.330 0.870 0.382 0.925 ;
      RECT 0.330 0.332 0.368 0.567 ;
      RECT 0.307 0.332 0.330 0.925 ;
      RECT 0.139 0.332 0.307 0.387 ;
      RECT 0.268 0.499 0.307 0.925 ;
      RECT 0.048 0.688 0.268 0.769 ;
      RECT 0.048 0.194 0.139 0.387 ;
  END
END ADDFX2

MACRO ADDFHX2
  CLASS CORE ;
  FOREIGN ADDFHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.900 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN S
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.797 0.219 5.845 0.494 ;
      RECT 5.797 0.627 5.812 0.958 ;
      RECT 5.755 0.219 5.797 0.958 ;
      RECT 5.737 0.357 5.755 0.958 ;
      RECT 5.723 0.654 5.737 0.958 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 5.466 0.331 5.514 0.412 ;
      RECT 5.424 0.331 5.466 0.761 ;
      RECT 5.406 0.344 5.424 0.761 ;
      RECT 5.262 0.706 5.406 0.761 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 4.994 0.546 5.169 0.649 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.588 0.635 3.699 0.715 ;
      RECT 3.527 0.635 3.588 0.761 ;
      RECT 3.363 0.635 3.527 0.715 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.191 0.433 0.327 0.571 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.655 -0.080 5.900 0.080 ;
      RECT 5.566 -0.080 5.655 0.211 ;
      RECT 5.314 -0.080 5.566 0.080 ;
      RECT 5.224 -0.080 5.314 0.122 ;
      RECT 3.570 -0.080 5.224 0.080 ;
      RECT 3.481 -0.080 3.570 0.122 ;
      RECT 0.881 -0.080 3.481 0.080 ;
      RECT 0.791 -0.080 0.881 0.122 ;
      RECT 0.350 -0.080 0.791 0.080 ;
      RECT 0.260 -0.080 0.350 0.122 ;
      RECT 0.000 -0.080 0.260 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.623 1.120 5.900 1.280 ;
      RECT 5.533 0.988 5.623 1.280 ;
      RECT 5.291 1.120 5.533 1.280 ;
      RECT 5.202 0.988 5.291 1.280 ;
      RECT 4.940 1.120 5.202 1.280 ;
      RECT 4.834 1.078 4.940 1.280 ;
      RECT 3.705 1.120 4.834 1.280 ;
      RECT 3.615 0.970 3.705 1.280 ;
      RECT 3.326 1.120 3.615 1.280 ;
      RECT 3.237 0.970 3.326 1.280 ;
      RECT 0.962 1.120 3.237 1.280 ;
      RECT 0.873 0.911 0.962 1.280 ;
      RECT 0.380 1.120 0.873 1.280 ;
      RECT 0.291 0.967 0.380 1.280 ;
      RECT 0.000 1.120 0.291 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.527 0.526 5.587 0.913 ;
      RECT 4.539 0.858 5.527 0.913 ;
      RECT 5.278 0.239 5.339 0.579 ;
      RECT 5.010 0.239 5.278 0.294 ;
      RECT 4.888 0.356 5.114 0.411 ;
      RECT 4.888 0.744 5.092 0.799 ;
      RECT 4.950 0.150 5.010 0.294 ;
      RECT 4.183 0.150 4.950 0.205 ;
      RECT 4.827 0.260 4.888 0.799 ;
      RECT 4.336 0.260 4.827 0.314 ;
      RECT 4.776 0.549 4.827 0.636 ;
      RECT 4.714 0.369 4.767 0.424 ;
      RECT 4.714 0.721 4.729 0.802 ;
      RECT 4.654 0.369 4.714 0.802 ;
      RECT 4.639 0.721 4.654 0.802 ;
      RECT 4.525 0.369 4.576 0.424 ;
      RECT 4.525 0.785 4.539 0.977 ;
      RECT 4.464 0.369 4.525 0.977 ;
      RECT 4.450 0.785 4.464 0.977 ;
      RECT 4.336 0.751 4.350 0.944 ;
      RECT 4.275 0.260 4.336 0.944 ;
      RECT 4.261 0.751 4.275 0.944 ;
      RECT 4.123 0.150 4.183 0.798 ;
      RECT 4.117 0.743 4.123 0.798 ;
      RECT 4.042 0.743 4.117 0.975 ;
      RECT 3.987 0.151 4.048 0.686 ;
      RECT 4.028 0.780 4.042 0.975 ;
      RECT 3.983 0.151 3.987 0.246 ;
      RECT 3.351 0.192 3.983 0.246 ;
      RECT 3.879 0.335 3.927 0.726 ;
      RECT 3.879 0.819 3.894 1.014 ;
      RECT 3.866 0.335 3.879 1.014 ;
      RECT 3.770 0.335 3.866 0.389 ;
      RECT 3.819 0.671 3.866 1.014 ;
      RECT 3.805 0.819 3.819 1.014 ;
      RECT 3.745 0.457 3.806 0.545 ;
      RECT 3.515 0.824 3.805 0.879 ;
      RECT 3.681 0.321 3.770 0.402 ;
      RECT 3.486 0.457 3.745 0.512 ;
      RECT 3.426 0.824 3.515 1.025 ;
      RECT 3.426 0.301 3.486 0.512 ;
      RECT 3.206 0.301 3.426 0.356 ;
      RECT 3.206 0.824 3.426 0.879 ;
      RECT 3.206 0.411 3.360 0.465 ;
      RECT 3.290 0.157 3.351 0.246 ;
      RECT 2.552 0.157 3.290 0.212 ;
      RECT 3.146 0.269 3.206 0.356 ;
      RECT 3.146 0.411 3.206 0.900 ;
      RECT 2.673 0.269 3.146 0.324 ;
      RECT 3.025 0.380 3.085 1.023 ;
      RECT 2.733 0.380 3.025 0.435 ;
      RECT 2.621 0.968 3.025 1.023 ;
      RECT 2.901 0.490 2.962 0.910 ;
      RECT 2.673 0.490 2.901 0.545 ;
      RECT 1.889 0.855 2.901 0.910 ;
      RECT 2.782 0.738 2.836 0.793 ;
      RECT 2.721 0.601 2.782 0.793 ;
      RECT 2.552 0.601 2.721 0.656 ;
      RECT 2.612 0.269 2.673 0.545 ;
      RECT 2.546 0.968 2.621 1.050 ;
      RECT 2.491 0.150 2.552 0.656 ;
      RECT 1.156 0.995 2.546 1.050 ;
      RECT 2.416 0.737 2.493 0.792 ;
      RECT 2.178 0.150 2.491 0.205 ;
      RECT 2.356 0.300 2.416 0.792 ;
      RECT 2.293 0.300 2.356 0.355 ;
      RECT 2.011 0.737 2.356 0.792 ;
      RECT 2.178 0.627 2.293 0.682 ;
      RECT 2.118 0.150 2.178 0.682 ;
      RECT 1.989 0.293 2.011 0.792 ;
      RECT 1.951 0.150 1.989 0.792 ;
      RECT 1.929 0.150 1.951 0.348 ;
      RECT 1.609 0.150 1.929 0.205 ;
      RECT 1.829 0.446 1.889 0.919 ;
      RECT 1.800 0.446 1.829 0.501 ;
      RECT 1.326 0.864 1.829 0.919 ;
      RECT 1.739 0.269 1.800 0.501 ;
      RECT 1.685 0.724 1.714 0.805 ;
      RECT 1.625 0.571 1.685 0.805 ;
      RECT 1.609 0.571 1.625 0.626 ;
      RECT 1.549 0.150 1.609 0.626 ;
      RECT 1.003 0.150 1.549 0.205 ;
      RECT 1.470 0.725 1.530 0.806 ;
      RECT 1.441 0.260 1.470 0.806 ;
      RECT 1.409 0.260 1.441 0.793 ;
      RECT 1.125 0.260 1.409 0.314 ;
      RECT 1.387 0.369 1.409 0.457 ;
      RECT 1.266 0.596 1.326 0.919 ;
      RECT 1.255 0.596 1.266 0.651 ;
      RECT 1.195 0.369 1.255 0.651 ;
      RECT 1.095 0.785 1.156 1.050 ;
      RECT 1.065 0.260 1.125 0.370 ;
      RECT 1.058 0.785 1.095 0.852 ;
      RECT 0.994 0.315 1.065 0.370 ;
      RECT 0.994 0.785 1.058 0.839 ;
      RECT 0.943 0.150 1.003 0.248 ;
      RECT 0.933 0.315 0.994 0.839 ;
      RECT 0.137 0.193 0.943 0.248 ;
      RECT 0.734 0.315 0.933 0.370 ;
      RECT 0.776 0.785 0.933 0.839 ;
      RECT 0.770 0.498 0.860 0.579 ;
      RECT 0.678 0.785 0.776 0.852 ;
      RECT 0.535 0.511 0.770 0.565 ;
      RECT 0.644 0.302 0.734 0.383 ;
      RECT 0.517 0.965 0.631 1.020 ;
      RECT 0.535 0.348 0.550 0.429 ;
      RECT 0.484 0.348 0.535 0.565 ;
      RECT 0.456 0.821 0.517 1.020 ;
      RECT 0.475 0.348 0.484 0.733 ;
      RECT 0.460 0.348 0.475 0.429 ;
      RECT 0.423 0.511 0.475 0.733 ;
      RECT 0.137 0.821 0.456 0.876 ;
      RECT 0.394 0.652 0.423 0.733 ;
      RECT 0.122 0.193 0.137 0.369 ;
      RECT 0.122 0.674 0.137 1.012 ;
      RECT 0.076 0.193 0.122 1.012 ;
      RECT 0.062 0.288 0.076 1.012 ;
      RECT 0.047 0.288 0.062 0.369 ;
      RECT 0.047 0.674 0.062 1.012 ;
  END
END ADDFHX2

MACRO MX3X2
  CLASS CORE ;
  FOREIGN MX3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.000 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN Y
  DIRECTION OUTPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.906 0.706 3.943 0.761 ;
      RECT 3.846 0.180 3.906 1.006 ;
      RECT 3.817 0.180 3.846 0.373 ;
      RECT 3.817 0.701 3.846 1.006 ;
     END
  END Y

  PIN S1
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 3.408 0.579 3.491 0.660 ;
      RECT 3.348 0.579 3.408 0.894 ;
      RECT 2.920 0.839 3.348 0.894 ;
      RECT 2.819 0.839 2.920 0.919 ;
     END
  END S1

  PIN S0
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.012 0.951 2.072 1.033 ;
      RECT 0.752 0.951 2.012 1.006 ;
      RECT 0.639 0.951 0.752 1.014 ;
      RECT 0.626 0.951 0.639 1.027 ;
      RECT 0.614 0.960 0.626 1.027 ;
      RECT 0.524 0.960 0.614 1.040 ;
     END
  END S0

  PIN C
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.111 0.433 0.200 0.550 ;
      RECT 0.037 0.433 0.111 0.549 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 1.570 0.433 1.702 0.540 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.437 0.525 2.572 0.633 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.701 -0.080 4.000 0.080 ;
      RECT 3.611 -0.080 3.701 0.210 ;
      RECT 2.592 -0.080 3.611 0.080 ;
      RECT 2.502 -0.080 2.592 0.122 ;
      RECT 1.599 -0.080 2.502 0.080 ;
      RECT 1.510 -0.080 1.599 0.122 ;
      RECT 1.138 -0.080 1.510 0.080 ;
      RECT 1.049 -0.080 1.138 0.122 ;
      RECT 0.137 -0.080 1.049 0.080 ;
      RECT 0.047 -0.080 0.137 0.364 ;
      RECT 0.000 -0.080 0.047 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.701 1.120 4.000 1.280 ;
      RECT 3.611 0.877 3.701 1.280 ;
      RECT 2.590 1.120 3.611 1.280 ;
      RECT 2.501 1.078 2.590 1.280 ;
      RECT 1.599 1.120 2.501 1.280 ;
      RECT 1.510 1.078 1.599 1.280 ;
      RECT 1.105 1.120 1.510 1.280 ;
      RECT 1.016 1.078 1.105 1.280 ;
      RECT 0.137 1.120 1.016 1.280 ;
      RECT 0.047 0.757 0.137 1.280 ;
      RECT 0.000 1.120 0.047 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.659 0.295 3.719 0.787 ;
      RECT 3.516 0.295 3.659 0.350 ;
      RECT 3.532 0.732 3.659 0.787 ;
      RECT 3.507 0.408 3.593 0.508 ;
      RECT 3.472 0.732 3.532 1.042 ;
      RECT 3.427 0.157 3.516 0.350 ;
      RECT 3.296 0.437 3.507 0.492 ;
      RECT 2.727 0.987 3.472 1.042 ;
      RECT 3.207 0.194 3.296 0.492 ;
      RECT 3.204 0.437 3.207 0.492 ;
      RECT 3.144 0.437 3.204 0.762 ;
      RECT 3.115 0.681 3.144 0.762 ;
      RECT 3.058 0.200 3.087 0.402 ;
      RECT 3.000 0.200 3.058 0.592 ;
      RECT 3.000 0.681 3.014 0.762 ;
      RECT 2.997 0.200 3.000 0.762 ;
      RECT 2.190 0.200 2.997 0.255 ;
      RECT 2.939 0.537 2.997 0.762 ;
      RECT 2.925 0.681 2.939 0.762 ;
      RECT 2.777 0.336 2.931 0.417 ;
      RECT 2.777 0.688 2.792 0.769 ;
      RECT 2.717 0.336 2.777 0.769 ;
      RECT 2.667 0.939 2.727 1.042 ;
      RECT 2.702 0.336 2.717 0.417 ;
      RECT 2.702 0.688 2.717 0.769 ;
      RECT 2.217 0.939 2.667 0.994 ;
      RECT 2.356 0.317 2.385 0.398 ;
      RECT 2.356 0.692 2.385 0.885 ;
      RECT 2.295 0.317 2.356 0.885 ;
      RECT 2.157 0.842 2.217 0.994 ;
      RECT 2.141 0.200 2.190 0.310 ;
      RECT 1.557 0.842 2.157 0.896 ;
      RECT 2.141 0.679 2.155 0.760 ;
      RECT 2.088 0.200 2.141 0.760 ;
      RECT 2.080 0.206 2.088 0.760 ;
      RECT 2.066 0.679 2.080 0.760 ;
      RECT 1.943 0.329 2.004 0.773 ;
      RECT 1.808 0.329 1.943 0.410 ;
      RECT 1.800 0.718 1.943 0.773 ;
      RECT 1.812 0.150 1.897 0.205 ;
      RECT 1.867 0.526 1.881 0.607 ;
      RECT 1.792 0.526 1.867 0.650 ;
      RECT 1.751 0.150 1.812 0.261 ;
      RECT 1.710 0.705 1.800 0.786 ;
      RECT 1.340 0.595 1.792 0.650 ;
      RECT 0.841 0.206 1.751 0.261 ;
      RECT 1.497 0.825 1.557 0.896 ;
      RECT 1.167 0.825 1.497 0.880 ;
      RECT 1.320 0.346 1.340 0.650 ;
      RECT 1.260 0.346 1.320 0.770 ;
      RECT 1.244 0.346 1.260 0.411 ;
      RECT 1.231 0.689 1.260 0.770 ;
      RECT 0.866 0.346 1.244 0.401 ;
      RECT 1.107 0.814 1.167 0.880 ;
      RECT 0.516 0.814 1.107 0.869 ;
      RECT 0.812 0.679 0.901 0.760 ;
      RECT 0.805 0.346 0.866 0.605 ;
      RECT 0.751 0.171 0.841 0.261 ;
      RECT 0.667 0.692 0.812 0.746 ;
      RECT 0.730 0.524 0.805 0.605 ;
      RECT 0.667 0.325 0.743 0.406 ;
      RECT 0.606 0.325 0.667 0.746 ;
      RECT 0.507 0.186 0.518 0.379 ;
      RECT 0.507 0.814 0.516 0.895 ;
      RECT 0.447 0.186 0.507 0.895 ;
      RECT 0.428 0.186 0.447 0.379 ;
      RECT 0.427 0.814 0.447 0.895 ;
      RECT 0.266 0.186 0.327 0.965 ;
      RECT 0.237 0.186 0.266 0.379 ;
      RECT 0.237 0.742 0.266 0.965 ;
  END
END MX3X2

MACRO TLATNTSCAX2
  CLASS CORE ;
  FOREIGN TLATNTSCAX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.300 BY 1.2 ;
  SYMMETRY X Y ;
  SITE CoreSite ;

  PIN ECK
  DIRECTION OUTPUT TRISTATE ;
     PORT
      LAYER Metal1 ;
      RECT 2.412 0.338 2.432 0.419 ;
      RECT 2.412 0.669 2.432 0.761 ;
      RECT 2.351 0.338 2.412 0.761 ;
      RECT 2.342 0.338 2.351 0.419 ;
      RECT 2.342 0.627 2.351 0.761 ;
      RECT 2.314 0.706 2.342 0.761 ;
     END
  END ECK

  PIN E
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 2.816 0.504 2.916 0.654 ;
     END
  END E

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
     PORT
      LAYER Metal1 ;
      RECT 2.992 0.433 3.089 0.580 ;
     END
  END CK

  PIN SE
  DIRECTION INPUT ;
     PORT
      LAYER Metal1 ;
      RECT 0.986 0.464 1.037 0.545 ;
      RECT 0.925 0.439 0.986 0.545 ;
      RECT 0.824 0.464 0.925 0.545 ;
     END
  END SE

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.026 -0.080 3.300 0.080 ;
      RECT 2.937 -0.080 3.026 0.122 ;
      RECT 2.042 -0.080 2.937 0.080 ;
      RECT 1.953 -0.080 2.042 0.122 ;
      RECT 1.618 -0.080 1.953 0.080 ;
      RECT 1.529 -0.080 1.618 0.122 ;
      RECT 0.976 -0.080 1.529 0.080 ;
      RECT 0.884 -0.080 0.976 0.200 ;
      RECT 0.347 -0.080 0.884 0.080 ;
      RECT 0.258 -0.080 0.347 0.122 ;
      RECT 0.000 -0.080 0.258 0.080 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.026 1.120 3.300 1.280 ;
      RECT 2.937 0.733 3.026 1.280 ;
      RECT 2.053 1.120 2.937 1.280 ;
      RECT 1.963 0.839 2.053 1.280 ;
      RECT 1.474 1.120 1.963 1.280 ;
      RECT 1.384 1.078 1.474 1.280 ;
      RECT 0.976 1.120 1.384 1.280 ;
      RECT 0.884 1.002 0.976 1.280 ;
      RECT 0.337 1.120 0.884 1.280 ;
      RECT 0.247 1.078 0.337 1.280 ;
      RECT 0.000 1.120 0.247 1.280 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.213 0.752 3.216 0.833 ;
      RECT 3.184 0.312 3.213 0.833 ;
      RECT 3.155 0.298 3.184 0.833 ;
      RECT 3.153 0.193 3.155 0.833 ;
      RECT 3.095 0.193 3.153 0.379 ;
      RECT 3.126 0.752 3.153 0.833 ;
      RECT 1.447 0.193 3.095 0.248 ;
      RECT 2.746 0.343 2.826 0.424 ;
      RECT 2.746 0.769 2.826 0.850 ;
      RECT 2.746 0.955 2.761 1.036 ;
      RECT 2.737 0.343 2.746 1.036 ;
      RECT 2.686 0.369 2.737 1.036 ;
      RECT 2.671 0.955 2.686 1.036 ;
      RECT 2.607 0.338 2.621 0.419 ;
      RECT 2.607 0.813 2.621 0.894 ;
      RECT 2.546 0.338 2.607 0.894 ;
      RECT 2.532 0.338 2.546 0.419 ;
      RECT 2.532 0.813 2.546 0.894 ;
      RECT 2.242 0.839 2.532 0.894 ;
      RECT 2.214 0.338 2.242 0.419 ;
      RECT 2.214 0.813 2.242 0.894 ;
      RECT 2.154 0.338 2.214 0.894 ;
      RECT 2.153 0.338 2.154 0.419 ;
      RECT 2.153 0.710 2.154 0.894 ;
      RECT 1.842 0.338 2.153 0.393 ;
      RECT 1.849 0.710 2.153 0.764 ;
      RECT 1.880 0.490 2.093 0.571 ;
      RECT 1.721 0.490 1.880 0.558 ;
      RECT 1.788 0.710 1.849 0.890 ;
      RECT 1.753 0.312 1.842 0.393 ;
      RECT 1.661 0.490 1.721 0.817 ;
      RECT 1.611 0.490 1.661 0.545 ;
      RECT 1.474 0.762 1.661 0.817 ;
      RECT 1.600 0.952 1.629 1.033 ;
      RECT 1.550 0.313 1.611 0.545 ;
      RECT 1.599 0.612 1.600 0.694 ;
      RECT 1.539 0.877 1.600 1.033 ;
      RECT 1.537 0.600 1.599 0.694 ;
      RECT 1.313 0.313 1.550 0.368 ;
      RECT 0.820 0.877 1.539 0.932 ;
      RECT 1.226 0.600 1.537 0.655 ;
      RECT 1.384 0.736 1.474 0.817 ;
      RECT 1.421 0.163 1.447 0.248 ;
      RECT 1.387 0.150 1.421 0.248 ;
      RECT 1.332 0.150 1.387 0.231 ;
      RECT 0.655 0.749 1.384 0.804 ;
      RECT 1.111 0.176 1.332 0.231 ;
      RECT 1.224 0.300 1.313 0.381 ;
      RECT 1.216 0.477 1.226 0.655 ;
      RECT 1.126 0.464 1.216 0.655 ;
      RECT 0.722 0.600 1.126 0.655 ;
      RECT 1.050 0.176 1.111 0.325 ;
      RECT 0.601 0.270 1.050 0.325 ;
      RECT 0.759 0.877 0.820 1.050 ;
      RECT 0.464 0.995 0.759 1.050 ;
      RECT 0.662 0.443 0.722 0.655 ;
      RECT 0.500 0.574 0.662 0.629 ;
      RECT 0.638 0.749 0.655 0.899 ;
      RECT 0.478 0.161 0.638 0.215 ;
      RECT 0.595 0.749 0.638 0.939 ;
      RECT 0.541 0.270 0.601 0.518 ;
      RECT 0.546 0.844 0.595 0.939 ;
      RECT 0.213 0.844 0.546 0.899 ;
      RECT 0.425 0.463 0.541 0.518 ;
      RECT 0.405 0.574 0.500 0.773 ;
      RECT 0.364 0.313 0.480 0.395 ;
      RECT 0.417 0.161 0.478 0.248 ;
      RECT 0.404 0.954 0.464 1.050 ;
      RECT 0.243 0.193 0.417 0.248 ;
      RECT 0.364 0.574 0.405 0.629 ;
      RECT 0.137 0.954 0.404 1.008 ;
      RECT 0.304 0.313 0.364 0.629 ;
      RECT 0.213 0.193 0.243 0.348 ;
      RECT 0.183 0.193 0.213 0.899 ;
      RECT 0.153 0.293 0.183 0.899 ;
      RECT 0.092 0.954 0.137 1.042 ;
      RECT 0.092 0.150 0.122 0.233 ;
      RECT 0.062 0.150 0.092 1.042 ;
      RECT 0.032 0.179 0.062 1.042 ;
  END
END TLATNTSCAX2

MACRO MEM1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM1 0 0 ;
  SIZE 426.965 BY 114.215 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal6 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal3 ;
        RECT 12.00 77.64 12.66 78.30 ;
      LAYER Metal4 ;
        RECT 12.00 77.64 12.66 78.30 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal6 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal3 ;
        RECT 12.00 71.52 12.66 72.18 ;
      LAYER Metal4 ;
        RECT 12.00 71.52 12.66 72.18 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal6 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal3 ;
        RECT 12.00 68.42 12.66 69.08 ;
      LAYER Metal4 ;
        RECT 12.00 68.42 12.66 69.08 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal6 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal3 ;
        RECT 12.00 62.30 12.66 62.96 ;
      LAYER Metal4 ;
        RECT 12.00 62.30 12.66 62.96 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal6 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal3 ;
        RECT 12.00 59.28 12.66 59.94 ;
      LAYER Metal4 ;
        RECT 12.00 59.28 12.66 59.94 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal6 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal3 ;
        RECT 12.00 56.18 12.66 56.84 ;
      LAYER Metal4 ;
        RECT 12.00 56.18 12.66 56.84 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal6 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal3 ;
        RECT 12.00 50.06 12.66 50.72 ;
      LAYER Metal4 ;
        RECT 12.00 50.06 12.66 50.72 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal6 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal3 ;
        RECT 12.00 47.04 12.66 47.70 ;
      LAYER Metal4 ;
        RECT 12.00 47.04 12.66 47.70 ;
    END
  END A[7]
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal6 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal3 ;
        RECT 228.44 12.00 229.09 12.66 ;
      LAYER Metal4 ;
        RECT 228.44 12.00 229.09 12.66 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal6 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal3 ;
        RECT 238.18 12.00 238.84 12.66 ;
      LAYER Metal4 ;
        RECT 238.18 12.00 238.84 12.66 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal6 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal3 ;
        RECT 20.48 12.00 21.14 12.66 ;
      LAYER Metal4 ;
        RECT 20.48 12.00 21.14 12.66 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal6 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal3 ;
        RECT 129.00 12.00 129.66 12.66 ;
      LAYER Metal4 ;
        RECT 129.00 12.00 129.66 12.66 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal6 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal3 ;
        RECT 137.04 12.00 137.70 12.66 ;
      LAYER Metal4 ;
        RECT 137.04 12.00 137.70 12.66 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal6 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal3 ;
        RECT 151.34 12.00 152.00 12.66 ;
      LAYER Metal4 ;
        RECT 151.34 12.00 152.00 12.66 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal6 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal3 ;
        RECT 159.38 12.00 160.04 12.66 ;
      LAYER Metal4 ;
        RECT 159.38 12.00 160.04 12.66 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal6 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal3 ;
        RECT 172.62 12.00 173.28 12.66 ;
      LAYER Metal4 ;
        RECT 172.62 12.00 173.28 12.66 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal6 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal3 ;
        RECT 180.66 12.00 181.32 12.66 ;
      LAYER Metal4 ;
        RECT 180.66 12.00 181.32 12.66 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal6 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal3 ;
        RECT 245.65 12.00 246.31 12.66 ;
      LAYER Metal4 ;
        RECT 245.65 12.00 246.31 12.66 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal6 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal3 ;
        RECT 253.69 12.00 254.34 12.66 ;
      LAYER Metal4 ;
        RECT 253.69 12.00 254.34 12.66 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal6 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal3 ;
        RECT 266.93 12.00 267.58 12.66 ;
      LAYER Metal4 ;
        RECT 266.93 12.00 267.58 12.66 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal6 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal3 ;
        RECT 274.96 12.00 275.62 12.66 ;
      LAYER Metal4 ;
        RECT 274.96 12.00 275.62 12.66 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal6 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal3 ;
        RECT 28.52 12.00 29.18 12.66 ;
      LAYER Metal4 ;
        RECT 28.52 12.00 29.18 12.66 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal6 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal3 ;
        RECT 289.26 12.00 289.93 12.66 ;
      LAYER Metal4 ;
        RECT 289.26 12.00 289.93 12.66 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal6 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal3 ;
        RECT 297.31 12.00 297.96 12.66 ;
      LAYER Metal4 ;
        RECT 297.31 12.00 297.96 12.66 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal6 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal3 ;
        RECT 310.55 12.00 311.20 12.66 ;
      LAYER Metal4 ;
        RECT 310.55 12.00 311.20 12.66 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal6 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal3 ;
        RECT 318.58 12.00 319.25 12.66 ;
      LAYER Metal4 ;
        RECT 318.58 12.00 319.25 12.66 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal6 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal3 ;
        RECT 332.88 12.00 333.55 12.66 ;
      LAYER Metal4 ;
        RECT 332.88 12.00 333.55 12.66 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal6 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal3 ;
        RECT 340.93 12.00 341.58 12.66 ;
      LAYER Metal4 ;
        RECT 340.93 12.00 341.58 12.66 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal6 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal3 ;
        RECT 354.17 12.00 354.82 12.66 ;
      LAYER Metal4 ;
        RECT 354.17 12.00 354.82 12.66 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal6 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal3 ;
        RECT 362.20 12.00 362.87 12.66 ;
      LAYER Metal4 ;
        RECT 362.20 12.00 362.87 12.66 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal6 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal3 ;
        RECT 376.50 12.00 377.17 12.66 ;
      LAYER Metal4 ;
        RECT 376.50 12.00 377.17 12.66 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal6 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal3 ;
        RECT 384.55 12.00 385.20 12.66 ;
      LAYER Metal4 ;
        RECT 384.55 12.00 385.20 12.66 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal6 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal3 ;
        RECT 41.76 12.00 42.42 12.66 ;
      LAYER Metal4 ;
        RECT 41.76 12.00 42.42 12.66 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal6 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal3 ;
        RECT 397.79 12.00 398.44 12.66 ;
      LAYER Metal4 ;
        RECT 397.79 12.00 398.44 12.66 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal6 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal3 ;
        RECT 405.82 12.00 406.49 12.66 ;
      LAYER Metal4 ;
        RECT 405.82 12.00 406.49 12.66 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal6 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal3 ;
        RECT 49.80 12.00 50.46 12.66 ;
      LAYER Metal4 ;
        RECT 49.80 12.00 50.46 12.66 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal6 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal3 ;
        RECT 64.10 12.00 64.76 12.66 ;
      LAYER Metal4 ;
        RECT 64.10 12.00 64.76 12.66 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal6 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal3 ;
        RECT 72.14 12.00 72.80 12.66 ;
      LAYER Metal4 ;
        RECT 72.14 12.00 72.80 12.66 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal6 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal3 ;
        RECT 85.38 12.00 86.04 12.66 ;
      LAYER Metal4 ;
        RECT 85.38 12.00 86.04 12.66 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal6 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal3 ;
        RECT 93.42 12.00 94.08 12.66 ;
      LAYER Metal4 ;
        RECT 93.42 12.00 94.08 12.66 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal6 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal3 ;
        RECT 107.72 12.00 108.38 12.66 ;
      LAYER Metal4 ;
        RECT 107.72 12.00 108.38 12.66 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal6 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal3 ;
        RECT 115.76 12.00 116.42 12.66 ;
      LAYER Metal4 ;
        RECT 115.76 12.00 116.42 12.66 ;
    END
  END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal6 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal3 ;
        RECT 23.06 12.00 23.72 12.66 ;
      LAYER Metal4 ;
        RECT 23.06 12.00 23.72 12.66 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal6 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal3 ;
        RECT 131.58 12.00 132.24 12.66 ;
      LAYER Metal4 ;
        RECT 131.58 12.00 132.24 12.66 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal6 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal3 ;
        RECT 134.46 12.00 135.12 12.66 ;
      LAYER Metal4 ;
        RECT 134.46 12.00 135.12 12.66 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal6 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal3 ;
        RECT 153.92 12.00 154.58 12.66 ;
      LAYER Metal4 ;
        RECT 153.92 12.00 154.58 12.66 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal6 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal3 ;
        RECT 156.80 12.00 157.46 12.66 ;
      LAYER Metal4 ;
        RECT 156.80 12.00 157.46 12.66 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal6 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal3 ;
        RECT 175.20 12.00 175.86 12.66 ;
      LAYER Metal4 ;
        RECT 175.20 12.00 175.86 12.66 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal6 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal3 ;
        RECT 178.08 12.00 178.74 12.66 ;
      LAYER Metal4 ;
        RECT 178.08 12.00 178.74 12.66 ;
    END
  END Q[15]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal6 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal3 ;
        RECT 248.22 12.00 248.88 12.66 ;
      LAYER Metal4 ;
        RECT 248.22 12.00 248.88 12.66 ;
    END
  END Q[16]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal6 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal3 ;
        RECT 251.10 12.00 251.76 12.66 ;
      LAYER Metal4 ;
        RECT 251.10 12.00 251.76 12.66 ;
    END
  END Q[17]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal6 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal3 ;
        RECT 269.50 12.00 270.17 12.66 ;
      LAYER Metal4 ;
        RECT 269.50 12.00 270.17 12.66 ;
    END
  END Q[18]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal6 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal3 ;
        RECT 272.38 12.00 273.05 12.66 ;
      LAYER Metal4 ;
        RECT 272.38 12.00 273.05 12.66 ;
    END
  END Q[19]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal6 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal3 ;
        RECT 25.94 12.00 26.60 12.66 ;
      LAYER Metal4 ;
        RECT 25.94 12.00 26.60 12.66 ;
    END
  END Q[1]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal6 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal3 ;
        RECT 291.85 12.00 292.50 12.66 ;
      LAYER Metal4 ;
        RECT 291.85 12.00 292.50 12.66 ;
    END
  END Q[20]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal6 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal3 ;
        RECT 294.73 12.00 295.38 12.66 ;
      LAYER Metal4 ;
        RECT 294.73 12.00 295.38 12.66 ;
    END
  END Q[21]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal6 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal3 ;
        RECT 313.12 12.00 313.79 12.66 ;
      LAYER Metal4 ;
        RECT 313.12 12.00 313.79 12.66 ;
    END
  END Q[22]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal6 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal3 ;
        RECT 316.00 12.00 316.67 12.66 ;
      LAYER Metal4 ;
        RECT 316.00 12.00 316.67 12.66 ;
    END
  END Q[23]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal6 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal3 ;
        RECT 335.46 12.00 336.12 12.66 ;
      LAYER Metal4 ;
        RECT 335.46 12.00 336.12 12.66 ;
    END
  END Q[24]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal6 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal3 ;
        RECT 338.35 12.00 339.00 12.66 ;
      LAYER Metal4 ;
        RECT 338.35 12.00 339.00 12.66 ;
    END
  END Q[25]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal6 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal3 ;
        RECT 356.75 12.00 357.40 12.66 ;
      LAYER Metal4 ;
        RECT 356.75 12.00 357.40 12.66 ;
    END
  END Q[26]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal6 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal3 ;
        RECT 359.62 12.00 360.29 12.66 ;
      LAYER Metal4 ;
        RECT 359.62 12.00 360.29 12.66 ;
    END
  END Q[27]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal6 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal3 ;
        RECT 379.08 12.00 379.75 12.66 ;
      LAYER Metal4 ;
        RECT 379.08 12.00 379.75 12.66 ;
    END
  END Q[28]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal6 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal3 ;
        RECT 381.96 12.00 382.62 12.66 ;
      LAYER Metal4 ;
        RECT 381.96 12.00 382.62 12.66 ;
    END
  END Q[29]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal6 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal3 ;
        RECT 44.34 12.00 45.00 12.66 ;
      LAYER Metal4 ;
        RECT 44.34 12.00 45.00 12.66 ;
    END
  END Q[2]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal6 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal3 ;
        RECT 400.37 12.00 401.02 12.66 ;
      LAYER Metal4 ;
        RECT 400.37 12.00 401.02 12.66 ;
    END
  END Q[30]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal6 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal3 ;
        RECT 403.25 12.00 403.90 12.66 ;
      LAYER Metal4 ;
        RECT 403.25 12.00 403.90 12.66 ;
    END
  END Q[31]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal6 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal3 ;
        RECT 47.22 12.00 47.88 12.66 ;
      LAYER Metal4 ;
        RECT 47.22 12.00 47.88 12.66 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal6 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal3 ;
        RECT 66.68 12.00 67.34 12.66 ;
      LAYER Metal4 ;
        RECT 66.68 12.00 67.34 12.66 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal6 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal3 ;
        RECT 69.56 12.00 70.22 12.66 ;
      LAYER Metal4 ;
        RECT 69.56 12.00 70.22 12.66 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal6 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal3 ;
        RECT 87.96 12.00 88.62 12.66 ;
      LAYER Metal4 ;
        RECT 87.96 12.00 88.62 12.66 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal6 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal3 ;
        RECT 90.84 12.00 91.50 12.66 ;
      LAYER Metal4 ;
        RECT 90.84 12.00 91.50 12.66 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal6 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal3 ;
        RECT 110.30 12.00 110.96 12.66 ;
      LAYER Metal4 ;
        RECT 110.30 12.00 110.96 12.66 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal6 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal3 ;
        RECT 113.18 12.00 113.84 12.66 ;
      LAYER Metal4 ;
        RECT 113.18 12.00 113.84 12.66 ;
    END
  END Q[9]
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal6 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal3 ;
        RECT 234.48 12.00 235.14 12.66 ;
      LAYER Metal4 ;
        RECT 234.48 12.00 235.14 12.66 ;
    END
  END WE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 109.22 426.96 114.22 ;
        RECT 0.00 0.00 426.96 5.00 ;
      LAYER Metal2 ;
        RECT 421.96 0.00 426.96 114.22 ;
        RECT 0.00 0.00 5.00 114.22 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 103.61 421.37 108.61 ;
        RECT 5.60 5.60 421.37 10.60 ;
      LAYER Metal2 ;
        RECT 416.37 5.60 421.37 108.61 ;
        RECT 5.60 5.60 10.60 108.61 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 415.01 102.02 ;
    LAYER Metal3 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal4 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal5 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
    LAYER Metal6 ;
#      RECT 12.00 12.00 415.01 102.02 ;
        RECT 12.84 12.84 415.01 102.02 ;
        RECT 12.00 12.00 20.30 46.86 ;
        RECT 21.32 12.00 22.88 102.02 ;
        RECT 23.90 12.00 25.76 102.02 ;
        RECT 26.78 12.00 28.34 102.02 ;
        RECT 29.36 12.00 41.58 102.02 ;
        RECT 42.60 12.00 44.16 102.02 ;
        RECT 45.18 12.00 47.04 102.02 ;
        RECT 48.06 12.00 49.62 102.02 ;
        RECT 50.64 12.00 63.92 102.02 ;
        RECT 64.94 12.00 66.50 102.02 ;
        RECT 67.52 12.00 69.38 102.02 ;
        RECT 70.40 12.00 71.96 102.02 ;
        RECT 72.98 12.00 85.20 102.02 ;
        RECT 86.22 12.00 87.78 102.02 ;
        RECT 88.80 12.00 90.66 102.02 ;
        RECT 91.68 12.00 93.24 102.02 ;
        RECT 94.26 12.00 107.54 102.02 ;
        RECT 108.56 12.00 110.12 102.02 ;
        RECT 111.14 12.00 113.00 102.02 ;
        RECT 114.02 12.00 115.58 102.02 ;
        RECT 116.60 12.00 128.82 102.02 ;
        RECT 129.84 12.00 131.40 102.02 ;
        RECT 132.42 12.00 134.28 102.02 ;
        RECT 135.30 12.00 136.86 102.02 ;
        RECT 137.88 12.00 151.16 102.02 ;
        RECT 152.18 12.00 153.74 102.02 ;
        RECT 154.76 12.00 156.62 102.02 ;
        RECT 157.64 12.00 159.20 102.02 ;
        RECT 160.22 12.00 172.44 102.02 ;
        RECT 173.46 12.00 175.02 102.02 ;
        RECT 176.04 12.00 177.90 102.02 ;
        RECT 178.92 12.00 180.48 102.02 ;
        RECT 181.50 12.00 228.26 102.02 ;
        RECT 229.27 12.00 234.30 102.02 ;
        RECT 235.32 12.00 238.00 102.02 ;
        RECT 239.02 12.00 245.47 102.02 ;
        RECT 246.49 12.00 248.04 102.02 ;
        RECT 249.06 12.00 250.92 102.02 ;
        RECT 251.94 12.00 253.51 102.02 ;
        RECT 254.52 12.00 266.75 102.02 ;
        RECT 267.76 12.00 269.32 102.02 ;
        RECT 270.35 12.00 272.20 102.02 ;
        RECT 273.23 12.00 274.78 102.02 ;
        RECT 275.80 12.00 289.08 102.02 ;
        RECT 290.11 12.00 291.67 102.02 ;
        RECT 292.68 12.00 294.55 102.02 ;
        RECT 295.56 12.00 297.13 102.02 ;
        RECT 298.14 12.00 310.37 102.02 ;
        RECT 311.38 12.00 312.94 102.02 ;
        RECT 313.97 12.00 315.82 102.02 ;
        RECT 316.85 12.00 318.40 102.02 ;
        RECT 319.43 12.00 332.70 102.02 ;
        RECT 333.73 12.00 335.28 102.02 ;
        RECT 336.30 12.00 338.17 102.02 ;
        RECT 339.18 12.00 340.75 102.02 ;
        RECT 341.76 12.00 353.99 102.02 ;
        RECT 355.00 12.00 356.57 102.02 ;
        RECT 357.58 12.00 359.44 102.02 ;
        RECT 360.47 12.00 362.02 102.02 ;
        RECT 363.05 12.00 376.32 102.02 ;
        RECT 377.35 12.00 378.90 102.02 ;
        RECT 379.93 12.00 381.78 102.02 ;
        RECT 382.80 12.00 384.37 102.02 ;
        RECT 385.38 12.00 397.61 102.02 ;
        RECT 398.62 12.00 400.19 102.02 ;
        RECT 401.20 12.00 403.07 102.02 ;
        RECT 404.08 12.00 405.64 102.02 ;
        RECT 406.67 12.00 415.01 102.02 ;
        RECT 12.00 47.88 415.01 49.88 ;
        RECT 12.00 50.90 415.01 56.00 ;
        RECT 12.00 57.02 415.01 59.10 ;
        RECT 12.00 60.12 415.01 62.12 ;
        RECT 12.00 63.14 415.01 68.24 ;
        RECT 12.00 69.26 415.01 71.34 ;
        RECT 12.00 72.36 415.01 77.46 ;
        RECT 12.00 78.48 415.01 102.02 ;
  END
END MEM1

MACRO MEM2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2 0 0 ;
  SIZE 423.015 BY 145.035 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal6 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal3 ;
        RECT 12.00 102.42 12.66 103.08 ;
      LAYER Metal4 ;
        RECT 12.00 102.42 12.66 103.08 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal6 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal3 ;
        RECT 12.00 96.30 12.66 96.96 ;
      LAYER Metal4 ;
        RECT 12.00 96.30 12.66 96.96 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal6 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal3 ;
        RECT 12.00 87.08 12.66 87.74 ;
      LAYER Metal4 ;
        RECT 12.00 87.08 12.66 87.74 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal6 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal3 ;
        RECT 12.00 84.06 12.66 84.72 ;
      LAYER Metal4 ;
        RECT 12.00 84.06 12.66 84.72 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal6 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal3 ;
        RECT 12.00 80.96 12.66 81.62 ;
      LAYER Metal4 ;
        RECT 12.00 80.96 12.66 81.62 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal6 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal3 ;
        RECT 12.00 74.84 12.66 75.50 ;
      LAYER Metal4 ;
        RECT 12.00 74.84 12.66 75.50 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal6 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal3 ;
        RECT 12.00 71.82 12.66 72.48 ;
      LAYER Metal4 ;
        RECT 12.00 71.82 12.66 72.48 ;
    END
  END A1[6]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal6 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal3 ;
        RECT 12.00 36.40 12.66 37.06 ;
      LAYER Metal4 ;
        RECT 12.00 36.40 12.66 37.06 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal6 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal3 ;
        RECT 12.00 42.52 12.66 43.18 ;
      LAYER Metal4 ;
        RECT 12.00 42.52 12.66 43.18 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal6 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal3 ;
        RECT 12.00 51.74 12.66 52.40 ;
      LAYER Metal4 ;
        RECT 12.00 51.74 12.66 52.40 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal6 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal3 ;
        RECT 12.00 54.76 12.66 55.42 ;
      LAYER Metal4 ;
        RECT 12.00 54.76 12.66 55.42 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal6 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal3 ;
        RECT 12.00 57.86 12.66 58.52 ;
      LAYER Metal4 ;
        RECT 12.00 57.86 12.66 58.52 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal6 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal3 ;
        RECT 12.00 63.98 12.66 64.64 ;
      LAYER Metal4 ;
        RECT 12.00 63.98 12.66 64.64 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal6 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal3 ;
        RECT 12.00 67.00 12.66 67.66 ;
      LAYER Metal4 ;
        RECT 12.00 67.00 12.66 67.66 ;
    END
  END A2[6]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal6 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal3 ;
        RECT 210.28 12.00 210.94 12.66 ;
      LAYER Metal4 ;
        RECT 210.28 12.00 210.94 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12.00 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12.00 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal6 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal3 ;
        RECT 218.91 12.00 219.56 12.66 ;
      LAYER Metal4 ;
        RECT 218.91 12.00 219.56 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal6 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal3 ;
        RECT 187.74 12.00 188.40 12.66 ;
      LAYER Metal4 ;
        RECT 187.74 12.00 188.40 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12.00 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12.00 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12.00 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12.00 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.40 12.00 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.40 12.00 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12.00 144.20 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12.00 144.20 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12.00 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12.00 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12.00 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12.00 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12.00 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12.00 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal6 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal3 ;
        RECT 221.68 12.00 222.34 12.66 ;
      LAYER Metal4 ;
        RECT 221.68 12.00 222.34 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal6 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal3 ;
        RECT 241.82 12.00 242.48 12.66 ;
      LAYER Metal4 ;
        RECT 241.82 12.00 242.48 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal6 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal3 ;
        RECT 242.96 12.00 243.62 12.66 ;
      LAYER Metal4 ;
        RECT 242.96 12.00 243.62 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal6 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal3 ;
        RECT 263.10 12.00 263.76 12.66 ;
      LAYER Metal4 ;
        RECT 263.10 12.00 263.76 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36.00 12.00 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36.00 12.00 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal6 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal3 ;
        RECT 264.24 12.00 264.90 12.66 ;
      LAYER Metal4 ;
        RECT 264.24 12.00 264.90 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal6 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal3 ;
        RECT 284.38 12.00 285.04 12.66 ;
      LAYER Metal4 ;
        RECT 284.38 12.00 285.04 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal6 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal3 ;
        RECT 285.52 12.00 286.18 12.66 ;
      LAYER Metal4 ;
        RECT 285.52 12.00 286.18 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal6 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal3 ;
        RECT 305.66 12.00 306.32 12.66 ;
      LAYER Metal4 ;
        RECT 305.66 12.00 306.32 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal6 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal3 ;
        RECT 306.80 12.00 307.46 12.66 ;
      LAYER Metal4 ;
        RECT 306.80 12.00 307.46 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal6 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal3 ;
        RECT 326.94 12.00 327.60 12.66 ;
      LAYER Metal4 ;
        RECT 326.94 12.00 327.60 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal6 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal3 ;
        RECT 328.08 12.00 328.74 12.66 ;
      LAYER Metal4 ;
        RECT 328.08 12.00 328.74 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal6 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal3 ;
        RECT 348.22 12.00 348.88 12.66 ;
      LAYER Metal4 ;
        RECT 348.22 12.00 348.88 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal6 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal3 ;
        RECT 349.36 12.00 350.02 12.66 ;
      LAYER Metal4 ;
        RECT 349.36 12.00 350.02 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal6 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal3 ;
        RECT 369.50 12.00 370.16 12.66 ;
      LAYER Metal4 ;
        RECT 369.50 12.00 370.16 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12.00 37.80 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12.00 37.80 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal6 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal3 ;
        RECT 370.64 12.00 371.30 12.66 ;
      LAYER Metal4 ;
        RECT 370.64 12.00 371.30 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal6 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal3 ;
        RECT 390.78 12.00 391.44 12.66 ;
      LAYER Metal4 ;
        RECT 390.78 12.00 391.44 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12.00 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12.00 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12.00 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12.00 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12.00 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12.00 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.70 12.00 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.70 12.00 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12.00 100.50 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12.00 100.50 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12.00 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12.00 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12.00 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12.00 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12.00 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12.00 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12.00 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12.00 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.90 12.00 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.90 12.00 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12.00 153.70 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12.00 153.70 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12.00 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12.00 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12.00 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12.00 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12.00 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12.00 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal6 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal3 ;
        RECT 231.18 12.00 231.84 12.66 ;
      LAYER Metal4 ;
        RECT 231.18 12.00 231.84 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal6 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal3 ;
        RECT 232.32 12.00 232.98 12.66 ;
      LAYER Metal4 ;
        RECT 232.32 12.00 232.98 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal6 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal3 ;
        RECT 252.46 12.00 253.12 12.66 ;
      LAYER Metal4 ;
        RECT 252.46 12.00 253.12 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal6 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal3 ;
        RECT 253.60 12.00 254.26 12.66 ;
      LAYER Metal4 ;
        RECT 253.60 12.00 254.26 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.50 12.00 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.50 12.00 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal6 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal3 ;
        RECT 273.74 12.00 274.40 12.66 ;
      LAYER Metal4 ;
        RECT 273.74 12.00 274.40 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal6 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal3 ;
        RECT 274.88 12.00 275.54 12.66 ;
      LAYER Metal4 ;
        RECT 274.88 12.00 275.54 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal6 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal3 ;
        RECT 295.02 12.00 295.68 12.66 ;
      LAYER Metal4 ;
        RECT 295.02 12.00 295.68 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal6 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal3 ;
        RECT 296.16 12.00 296.82 12.66 ;
      LAYER Metal4 ;
        RECT 296.16 12.00 296.82 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal6 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal3 ;
        RECT 316.30 12.00 316.96 12.66 ;
      LAYER Metal4 ;
        RECT 316.30 12.00 316.96 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal6 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal3 ;
        RECT 317.44 12.00 318.10 12.66 ;
      LAYER Metal4 ;
        RECT 317.44 12.00 318.10 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal6 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal3 ;
        RECT 337.58 12.00 338.24 12.66 ;
      LAYER Metal4 ;
        RECT 337.58 12.00 338.24 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal6 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal3 ;
        RECT 338.72 12.00 339.38 12.66 ;
      LAYER Metal4 ;
        RECT 338.72 12.00 339.38 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal6 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal3 ;
        RECT 358.86 12.00 359.52 12.66 ;
      LAYER Metal4 ;
        RECT 358.86 12.00 359.52 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal6 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal3 ;
        RECT 360.00 12.00 360.66 12.66 ;
      LAYER Metal4 ;
        RECT 360.00 12.00 360.66 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12.00 47.30 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12.00 47.30 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal6 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal3 ;
        RECT 380.14 12.00 380.80 12.66 ;
      LAYER Metal4 ;
        RECT 380.14 12.00 380.80 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal6 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal3 ;
        RECT 381.28 12.00 381.94 12.66 ;
      LAYER Metal4 ;
        RECT 381.28 12.00 381.94 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12.00 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12.00 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12.00 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12.00 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12.00 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12.00 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.20 12.00 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.20 12.00 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12.00 91.00 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12.00 91.00 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12.00 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12.00 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12.00 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12.00 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12.00 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12.00 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12.00 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12.00 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.10 12.00 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.10 12.00 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12.00 147.50 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12.00 147.50 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12.00 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12.00 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12.00 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12.00 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12.00 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12.00 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal6 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal3 ;
        RECT 224.98 12.00 225.64 12.66 ;
      LAYER Metal4 ;
        RECT 224.98 12.00 225.64 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal6 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal3 ;
        RECT 238.52 12.00 239.18 12.66 ;
      LAYER Metal4 ;
        RECT 238.52 12.00 239.18 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal6 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal3 ;
        RECT 246.26 12.00 246.92 12.66 ;
      LAYER Metal4 ;
        RECT 246.26 12.00 246.92 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal6 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal3 ;
        RECT 259.80 12.00 260.46 12.66 ;
      LAYER Metal4 ;
        RECT 259.80 12.00 260.46 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.70 12.00 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.70 12.00 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal6 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal3 ;
        RECT 267.54 12.00 268.20 12.66 ;
      LAYER Metal4 ;
        RECT 267.54 12.00 268.20 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal6 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal3 ;
        RECT 281.08 12.00 281.74 12.66 ;
      LAYER Metal4 ;
        RECT 281.08 12.00 281.74 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal6 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal3 ;
        RECT 288.82 12.00 289.48 12.66 ;
      LAYER Metal4 ;
        RECT 288.82 12.00 289.48 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal6 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal3 ;
        RECT 302.36 12.00 303.02 12.66 ;
      LAYER Metal4 ;
        RECT 302.36 12.00 303.02 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal6 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal3 ;
        RECT 310.10 12.00 310.76 12.66 ;
      LAYER Metal4 ;
        RECT 310.10 12.00 310.76 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal6 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal3 ;
        RECT 323.64 12.00 324.30 12.66 ;
      LAYER Metal4 ;
        RECT 323.64 12.00 324.30 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal6 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal3 ;
        RECT 331.38 12.00 332.04 12.66 ;
      LAYER Metal4 ;
        RECT 331.38 12.00 332.04 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal6 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal3 ;
        RECT 344.92 12.00 345.58 12.66 ;
      LAYER Metal4 ;
        RECT 344.92 12.00 345.58 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal6 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal3 ;
        RECT 352.66 12.00 353.32 12.66 ;
      LAYER Metal4 ;
        RECT 352.66 12.00 353.32 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal6 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal3 ;
        RECT 366.20 12.00 366.86 12.66 ;
      LAYER Metal4 ;
        RECT 366.20 12.00 366.86 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12.00 41.10 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12.00 41.10 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal6 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal3 ;
        RECT 373.94 12.00 374.60 12.66 ;
      LAYER Metal4 ;
        RECT 373.94 12.00 374.60 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal6 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal3 ;
        RECT 388.36 12.00 389.02 12.66 ;
      LAYER Metal4 ;
        RECT 388.36 12.00 389.02 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12.00 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12.00 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12.00 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12.00 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12.00 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12.00 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83.00 12.00 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83.00 12.00 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12.00 97.20 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12.00 97.20 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12.00 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12.00 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12.00 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12.00 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12.00 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12.00 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12.00 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12.00 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.20 12.00 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.20 12.00 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12.00 150.40 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12.00 150.40 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12.00 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12.00 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12.00 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12.00 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12.00 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12.00 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal6 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal3 ;
        RECT 227.88 12.00 228.54 12.66 ;
      LAYER Metal4 ;
        RECT 227.88 12.00 228.54 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal6 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal3 ;
        RECT 235.62 12.00 236.28 12.66 ;
      LAYER Metal4 ;
        RECT 235.62 12.00 236.28 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal6 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal3 ;
        RECT 249.16 12.00 249.82 12.66 ;
      LAYER Metal4 ;
        RECT 249.16 12.00 249.82 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal6 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal3 ;
        RECT 256.90 12.00 257.56 12.66 ;
      LAYER Metal4 ;
        RECT 256.90 12.00 257.56 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.80 12.00 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.80 12.00 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal6 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal3 ;
        RECT 270.44 12.00 271.10 12.66 ;
      LAYER Metal4 ;
        RECT 270.44 12.00 271.10 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal6 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal3 ;
        RECT 278.18 12.00 278.84 12.66 ;
      LAYER Metal4 ;
        RECT 278.18 12.00 278.84 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal6 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal3 ;
        RECT 291.72 12.00 292.38 12.66 ;
      LAYER Metal4 ;
        RECT 291.72 12.00 292.38 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal6 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal3 ;
        RECT 299.46 12.00 300.12 12.66 ;
      LAYER Metal4 ;
        RECT 299.46 12.00 300.12 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal6 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal3 ;
        RECT 313.00 12.00 313.66 12.66 ;
      LAYER Metal4 ;
        RECT 313.00 12.00 313.66 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal6 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal3 ;
        RECT 320.74 12.00 321.40 12.66 ;
      LAYER Metal4 ;
        RECT 320.74 12.00 321.40 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal6 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal3 ;
        RECT 334.28 12.00 334.94 12.66 ;
      LAYER Metal4 ;
        RECT 334.28 12.00 334.94 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal6 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal3 ;
        RECT 342.02 12.00 342.68 12.66 ;
      LAYER Metal4 ;
        RECT 342.02 12.00 342.68 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal6 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal3 ;
        RECT 355.56 12.00 356.22 12.66 ;
      LAYER Metal4 ;
        RECT 355.56 12.00 356.22 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal6 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal3 ;
        RECT 363.30 12.00 363.96 12.66 ;
      LAYER Metal4 ;
        RECT 363.30 12.00 363.96 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12.00 44.00 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12.00 44.00 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal6 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal3 ;
        RECT 376.84 12.00 377.50 12.66 ;
      LAYER Metal4 ;
        RECT 376.84 12.00 377.50 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal6 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal3 ;
        RECT 384.58 12.00 385.24 12.66 ;
      LAYER Metal4 ;
        RECT 384.58 12.00 385.24 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12.00 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12.00 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12.00 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12.00 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12.00 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12.00 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.90 12.00 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.90 12.00 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12.00 94.30 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12.00 94.30 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12.00 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12.00 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12.00 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12.00 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal6 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal3 ;
        RECT 212.68 12.00 213.34 12.66 ;
      LAYER Metal4 ;
        RECT 212.68 12.00 213.34 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12.00 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12.00 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0.00 140.03 423.01 145.03 ;
        RECT 0.00 0.00 423.01 5.00 ;
      LAYER Metal2 ;
        RECT 418.01 0.00 423.01 145.03 ;
        RECT 0.00 0.00 5.00 145.03 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.60 134.44 417.42 139.44 ;
        RECT 5.60 5.60 417.42 10.60 ;
      LAYER Metal2 ;
        RECT 412.42 5.60 417.42 139.44 ;
        RECT 5.60 5.60 10.60 139.44 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal2 ;
      RECT 12.00 12.00 411.02 132.97 ;
    LAYER Metal3 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal4 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal5 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
    LAYER Metal6 ;
#      RECT 12.00 12.00 411.02 132.97 ;
        RECT 12.84 12.84 411.02 132.97 ;
        RECT 12.00 12.00 15.68 36.22 ;
        RECT 16.70 12.00 18.10 132.97 ;
        RECT 19.12 12.00 21.88 132.97 ;
        RECT 22.90 12.00 25.18 132.97 ;
        RECT 26.20 12.00 26.32 132.97 ;
        RECT 27.34 12.00 29.62 132.97 ;
        RECT 30.64 12.00 32.52 132.97 ;
        RECT 33.54 12.00 35.82 132.97 ;
        RECT 36.84 12.00 36.96 132.97 ;
        RECT 37.98 12.00 40.26 132.97 ;
        RECT 41.28 12.00 43.16 132.97 ;
        RECT 44.18 12.00 46.46 132.97 ;
        RECT 47.48 12.00 47.60 132.97 ;
        RECT 48.62 12.00 50.90 132.97 ;
        RECT 51.92 12.00 53.80 132.97 ;
        RECT 54.82 12.00 57.10 132.97 ;
        RECT 58.12 12.00 58.24 132.97 ;
        RECT 59.26 12.00 61.54 132.97 ;
        RECT 62.56 12.00 64.44 132.97 ;
        RECT 65.46 12.00 67.74 132.97 ;
        RECT 68.76 12.00 68.88 132.97 ;
        RECT 69.90 12.00 72.18 132.97 ;
        RECT 73.20 12.00 75.08 132.97 ;
        RECT 76.10 12.00 78.38 132.97 ;
        RECT 79.40 12.00 79.52 132.97 ;
        RECT 80.54 12.00 82.82 132.97 ;
        RECT 83.84 12.00 85.72 132.97 ;
        RECT 86.74 12.00 89.02 132.97 ;
        RECT 90.04 12.00 90.16 132.97 ;
        RECT 91.18 12.00 93.46 132.97 ;
        RECT 94.48 12.00 96.36 132.97 ;
        RECT 97.38 12.00 99.66 132.97 ;
        RECT 100.68 12.00 100.80 132.97 ;
        RECT 101.82 12.00 104.10 132.97 ;
        RECT 105.12 12.00 107.00 132.97 ;
        RECT 108.02 12.00 110.30 132.97 ;
        RECT 111.32 12.00 111.44 132.97 ;
        RECT 112.46 12.00 114.74 132.97 ;
        RECT 115.76 12.00 117.64 132.97 ;
        RECT 118.66 12.00 120.94 132.97 ;
        RECT 121.96 12.00 122.08 132.97 ;
        RECT 123.10 12.00 125.38 132.97 ;
        RECT 126.40 12.00 128.28 132.97 ;
        RECT 129.30 12.00 131.58 132.97 ;
        RECT 132.60 12.00 132.72 132.97 ;
        RECT 133.74 12.00 136.02 132.97 ;
        RECT 137.04 12.00 138.92 132.97 ;
        RECT 139.94 12.00 142.22 132.97 ;
        RECT 143.24 12.00 143.36 132.97 ;
        RECT 144.38 12.00 146.66 132.97 ;
        RECT 147.68 12.00 149.56 132.97 ;
        RECT 150.58 12.00 152.86 132.97 ;
        RECT 153.88 12.00 154.00 132.97 ;
        RECT 155.02 12.00 157.30 132.97 ;
        RECT 158.32 12.00 160.20 132.97 ;
        RECT 161.22 12.00 163.50 132.97 ;
        RECT 164.52 12.00 164.64 132.97 ;
        RECT 165.66 12.00 167.94 132.97 ;
        RECT 168.96 12.00 170.84 132.97 ;
        RECT 171.86 12.00 174.14 132.97 ;
        RECT 175.16 12.00 175.28 132.97 ;
        RECT 176.30 12.00 178.58 132.97 ;
        RECT 179.60 12.00 181.48 132.97 ;
        RECT 182.50 12.00 184.78 132.97 ;
        RECT 185.80 12.00 187.56 132.97 ;
        RECT 188.58 12.00 193.78 132.97 ;
        RECT 194.80 12.00 196.18 132.97 ;
        RECT 197.20 12.00 210.10 132.97 ;
        RECT 211.12 12.00 212.50 132.97 ;
        RECT 213.52 12.00 218.73 132.97 ;
        RECT 219.74 12.00 221.50 132.97 ;
        RECT 222.52 12.00 224.80 132.97 ;
        RECT 225.82 12.00 227.70 132.97 ;
        RECT 228.72 12.00 231.00 132.97 ;
        RECT 232.02 12.00 232.14 132.97 ;
        RECT 233.16 12.00 235.44 132.97 ;
        RECT 236.46 12.00 238.34 132.97 ;
        RECT 239.36 12.00 241.64 132.97 ;
        RECT 242.66 12.00 242.78 132.97 ;
        RECT 243.80 12.00 246.08 132.97 ;
        RECT 247.10 12.00 248.98 132.97 ;
        RECT 250.00 12.00 252.28 132.97 ;
        RECT 253.30 12.00 253.42 132.97 ;
        RECT 254.44 12.00 256.72 132.97 ;
        RECT 257.74 12.00 259.62 132.97 ;
        RECT 260.64 12.00 262.92 132.97 ;
        RECT 263.94 12.00 264.06 132.97 ;
        RECT 265.08 12.00 267.36 132.97 ;
        RECT 268.38 12.00 270.26 132.97 ;
        RECT 271.28 12.00 273.56 132.97 ;
        RECT 274.58 12.00 274.70 132.97 ;
        RECT 275.72 12.00 278.00 132.97 ;
        RECT 279.02 12.00 280.90 132.97 ;
        RECT 281.92 12.00 284.20 132.97 ;
        RECT 285.22 12.00 285.34 132.97 ;
        RECT 286.36 12.00 288.64 132.97 ;
        RECT 289.66 12.00 291.54 132.97 ;
        RECT 292.56 12.00 294.84 132.97 ;
        RECT 295.86 12.00 295.98 132.97 ;
        RECT 297.00 12.00 299.28 132.97 ;
        RECT 300.30 12.00 302.18 132.97 ;
        RECT 303.20 12.00 305.48 132.97 ;
        RECT 306.50 12.00 306.62 132.97 ;
        RECT 307.64 12.00 309.92 132.97 ;
        RECT 310.94 12.00 312.82 132.97 ;
        RECT 313.84 12.00 316.12 132.97 ;
        RECT 317.14 12.00 317.26 132.97 ;
        RECT 318.28 12.00 320.56 132.97 ;
        RECT 321.58 12.00 323.46 132.97 ;
        RECT 324.48 12.00 326.76 132.97 ;
        RECT 327.78 12.00 327.90 132.97 ;
        RECT 328.92 12.00 331.20 132.97 ;
        RECT 332.22 12.00 334.10 132.97 ;
        RECT 335.12 12.00 337.40 132.97 ;
        RECT 338.42 12.00 338.54 132.97 ;
        RECT 339.56 12.00 341.84 132.97 ;
        RECT 342.86 12.00 344.74 132.97 ;
        RECT 345.76 12.00 348.04 132.97 ;
        RECT 349.06 12.00 349.18 132.97 ;
        RECT 350.20 12.00 352.48 132.97 ;
        RECT 353.50 12.00 355.38 132.97 ;
        RECT 356.40 12.00 358.68 132.97 ;
        RECT 359.70 12.00 359.82 132.97 ;
        RECT 360.84 12.00 363.12 132.97 ;
        RECT 364.14 12.00 366.02 132.97 ;
        RECT 367.04 12.00 369.32 132.97 ;
        RECT 370.34 12.00 370.46 132.97 ;
        RECT 371.48 12.00 373.76 132.97 ;
        RECT 374.78 12.00 376.66 132.97 ;
        RECT 377.68 12.00 379.96 132.97 ;
        RECT 380.98 12.00 381.10 132.97 ;
        RECT 382.12 12.00 384.40 132.97 ;
        RECT 385.42 12.00 388.18 132.97 ;
        RECT 389.20 12.00 390.60 132.97 ;
        RECT 391.62 12.00 411.02 132.97 ;
        RECT 12.00 37.24 411.02 42.34 ;
        RECT 12.00 43.36 411.02 51.56 ;
        RECT 12.00 52.58 411.02 54.58 ;
        RECT 12.00 55.60 411.02 57.68 ;
        RECT 12.00 58.70 411.02 63.80 ;
        RECT 12.00 64.82 411.02 66.82 ;
        RECT 12.00 67.84 411.02 71.64 ;
        RECT 12.00 72.66 411.02 74.66 ;
        RECT 12.00 75.68 411.02 80.78 ;
        RECT 12.00 81.80 411.02 83.88 ;
        RECT 12.00 84.90 411.02 86.90 ;
        RECT 12.00 87.92 411.02 96.12 ;
        RECT 12.00 97.14 411.02 102.24 ;
        RECT 12.00 103.26 411.02 132.97 ;
  END
END MEM2

END LIBRARY

